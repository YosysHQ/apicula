`define PLL_DEVICE "GW1N-1"
`define PLL_FCLKIN "24"
`define PLL_FBDIV_SEL 9
`define PLL_IDIV_SEL  2
`define PLL_ODIV_SEL  8

