`define PLL_DEVICE "GW1N-1"
`define PLL_FCLKIN "24"
`define PLL_FBDIV_SEL 12
`define PLL_IDIV_SEL  5
`define PLL_ODIV_SEL  8

