`define PLL_DYN
`define PLL_DEVICE "GW1NSR-4C"
`define PLL_FCLKIN "12"
`define PLL_ODIV_SEL  64

`define PLL_FBDIV_SEL 12
`define PLL_IDIV_SEL  5

`define PLL_FBDIV_SEL_1 9
`define PLL_IDIV_SEL_1  2

// LCD
`define PLL_FBDIV_SEL_LCD 1
`define PLL_IDIV_SEL_LCD  2
