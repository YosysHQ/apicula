`define PLL_FCLKIN "50"

// LCD
`define PLL_FBDIV_SEL_LCD	1
`define PLL_ODIV0_SEL		32  // 25.2 MHz
`define PLL_IDIV_SEL_LCD	1

