../img-rom.vh