../img-video-ram1.vh