module top(R1C32_IOA);
inout R1C32_IOA;
wire R6C16_GBO1;
wire R8C38_GB10;
wire R4C6_GB00;
wire R27C26_GB70;
wire R10C34_W81;
wire R1C28_S26;
wire R15C42_GB60;
wire R10C29_CLK1;
wire R14C28_GB30;
wire R28C4_E81;
wire R7C46_GT10;
wire R13C19_GT00;
wire R14C2_GB20;
wire R1C1_C3;
wire R22C27_GB00;
wire R25C3_GB60;
wire R24C2_GB00;
wire R4C35_GB10;
wire R28C22_W10;
wire R6C10_GBO0;
wire R8C23_GT10;
wire R10C19_E83;
wire R12C11_GB60;
wire R27C15_GBO0;
wire R16C41_GB20;
wire R15C28_GT10;
wire R28C46_X06;
wire R9C37_GBO1;
wire R13C31_GB20;
wire R17C43_GB60;
wire R8C12_GB40;
wire R6C9_GBO0;
wire R25C20_GBO0;
wire R13C27_GBO1;
wire R1C47_CE2;
wire R10C25_F2;
wire R10C13_Q7;
wire R23C23_GB10;
wire R6C40_GBO1;
wire R7C25_GB30;
wire R16C6_GB10;
wire R10C13_CLK1;
wire R11C40_GB70;
wire R21C40_GB00;
wire R16C17_GB40;
wire R28C25_D4;
wire R13C46_GT00;
wire R23C6_GB70;
wire R11C23_GB30;
wire R9C11_GT00;
wire R24C16_GT00;
wire R22C29_GT10;
wire R9C2_GB50;
wire R6C7_GBO0;
wire R10C34_S11;
wire R25C26_GT10;
wire R11C37_GB50;
wire R28C19_C0;
wire R28C10_X02;
wire R28C40_W82;
wire R10C25_D3;
wire R1C47_W10;
wire R23C12_GB00;
wire R17C41_GB50;
wire R28C37_D5;
wire R28C22_Q7;
wire R9C4_GB20;
wire R3C8_GB20;
wire R25C24_GB30;
wire R21C33_GB20;
wire R28C37_EW20;
wire R14C13_GT00;
wire R7C39_GB30;
wire R4C44_GT00;
wire R10C25_S22;
wire R10C16_S23;
wire R10C16_X05;
wire R23C6_GBO1;
wire R16C31_GB30;
wire R28C7_S81;
wire R9C10_GB70;
wire R3C40_GB00;
wire R28C25_A5;
wire R10C25_F5;
wire R18C40_GBO0;
wire R23C16_GBO1;
wire R10C7_S24;
wire R2C9_GB00;
wire R10C22_A4;
wire R22C40_GB50;
wire R17C41_GT00;
wire R13C20_GB10;
wire R26C16_GB60;
wire R29C28_E82;
wire R13C43_GBO1;
wire R10C31_W20;
wire R28C37_B0;
wire R15C24_GB10;
wire R13C11_GBO0;
wire R11C2_GB20;
wire R24C14_GB40;
wire R4C26_GBO1;
wire R13C18_GB10;
wire R12C17_GBO1;
wire R15C4_GB70;
wire R28C10_B4;
wire R3C17_GB10;
wire R21C26_GB20;
wire R5C38_GB70;
wire R23C25_GBO1;
wire R3C36_GT00;
wire R24C2_GB60;
wire R8C15_GB30;
wire R21C12_GB10;
wire R10C34_N10;
wire R11C31_GB20;
wire R3C28_GB70;
wire R21C22_GB40;
wire R18C22_GT10;
wire R28C10_D0;
wire R22C20_GBO1;
wire R16C25_GBO1;
wire R24C8_GT00;
wire R25C27_GBO0;
wire R11C25_GBO1;
wire R1C32_S11;
wire R10C40_N23;
wire R24C13_GT10;
wire R12C40_GT00;
wire R8C46_GB10;
wire R9C46_GB30;
wire R5C43_GB60;
wire R18C11_GB70;
wire R11C44_GB10;
wire R3C25_GB70;
wire R10C37_E13;
wire R3C27_GB40;
wire R10C37_C1;
wire R16C11_GT10;
wire R26C17_GBO0;
wire R5C22_GB30;
wire R15C31_GT00;
wire R20C32_GT10;
wire R2C7_GBO0;
wire R6C39_GB60;
wire R4C39_GT00;
wire R6C37_GBO1;
wire R23C40_GBO1;
wire R10C34_Q2;
wire R7C7_GB10;
wire R17C30_GB60;
wire R28C46_Q0;
wire R28C37_F7;
wire R14C25_GB00;
wire R6C25_GT00;
wire R2C4_GB70;
wire R1C28_B6;
wire R23C26_GB50;
wire R17C33_GB10;
wire R7C14_GBO0;
wire R18C8_GB50;
wire R21C19_GT10;
wire R2C21_SPINE11;
wire R22C26_GB60;
wire R10C26_A1;
wire R24C41_GT10;
wire R24C36_GBO0;
wire R27C44_GBO1;
wire R26C17_GT00;
wire R18C9_GB10;
wire R20C11_GT00;
wire R21C26_GB30;
wire R26C20_GT00;
wire R17C21_GBO1;
wire R18C6_GB60;
wire R28C25_S26;
wire R7C21_GB50;
wire R5C31_GB20;
wire R14C28_GB20;
wire R7C34_GB10;
wire R1C32_W26;
wire R10C25_E12;
wire R9C45_GT10;
wire R28C34_CLK1;
wire R8C15_GBO0;
wire R10C25_A0;
wire R28C40_N11;
wire R21C30_GBO0;
wire R14C6_GB10;
wire R25C32_GB00;
wire R1C28_W26;
wire R28C16_Q5;
wire R8C5_GT00;
wire R6C21_GB60;
wire R27C38_GB50;
wire R11C11_GB10;
wire R18C26_GBO0;
wire R21C39_GT00;
wire R20C15_SPINE21;
wire R12C21_GB60;
wire R27C12_GB50;
wire R21C14_GB60;
wire R2C32_GB40;
wire R7C42_GB40;
wire R20C45_GT10;
wire R4C12_GB30;
wire R11C8_GB30;
wire R5C41_GB40;
wire R27C27_GB40;
wire R14C15_GT10;
wire R28C46_N24;
wire R4C3_GBO1;
wire R8C23_GB60;
wire R6C18_GT00;
wire R13C19_GBO1;
wire R22C21_GB70;
wire R16C43_GB60;
wire R29C28_SEL3;
wire R25C17_GB10;
wire R22C35_GB30;
wire R16C18_GT00;
wire R21C27_GT10;
wire R9C12_GB40;
wire R4C37_GB30;
wire R14C8_GBO0;
wire R1C32_F3;
wire R28C28_A4;
wire R28C34_A1;
wire R4C10_GB40;
wire R28C43_N22;
wire R28C7_S27;
wire R10C40_D5;
wire R15C22_GB30;
wire R24C24_GB60;
wire R15C36_GB50;
wire R10C26_N11;
wire R28C13_W11;
wire R25C24_GBO1;
wire R15C35_GB40;
wire R12C29_GT00;
wire R24C42_GB00;
wire R12C33_GT00;
wire R10C37_F6;
wire R8C21_GT00;
wire R14C4_GB10;
wire R11C14_GB00;
wire R16C29_GBO1;
wire R28C28_E80;
wire R28C31_D5;
wire R16C39_GB50;
wire R15C13_GB30;
wire R10C19_N23;
wire R10C13_C6;
wire R17C32_GB60;
wire R28C7_B0;
wire R13C3_GB20;
wire R14C37_GT00;
wire R13C3_GB60;
wire R10C22_C2;
wire R11C39_GB60;
wire R14C4_GBO1;
wire R28C28_E20;
wire R16C9_GT00;
wire R7C12_GBO0;
wire R7C7_GB40;
wire R10C30_N80;
wire R4C29_GB50;
wire R20C46_GBO1;
wire R10C31_A0;
wire R7C21_GT00;
wire R26C32_GT10;
wire R10C26_E12;
wire R28C7_N81;
wire R10C28_CLK0;
wire R2C9_GB50;
wire R28C7_D4;
wire R12C22_GT00;
wire R9C41_GT10;
wire R10C29_UNK127;
wire R7C7_GB20;
wire R5C32_GT00;
wire R18C23_GBO0;
wire R18C40_GBO1;
wire R2C18_GB00;
wire R26C12_GB60;
wire R10C13_SEL4;
wire R6C28_GB00;
wire R10C13_W13;
wire R18C45_GBO1;
wire R8C22_GB10;
wire R2C21_GB50;
wire R5C45_GB50;
wire R28C10_N20;
wire R10C29_A2;
wire R7C12_GT10;
wire R1C28_A2;
wire R3C33_GT00;
wire R26C8_GB20;
wire R2C6_GT10;
wire R28C22_SEL2;
wire R20C15_GBO0;
wire R18C14_GB40;
wire R22C13_GB50;
wire R25C18_GB60;
wire R12C34_GB70;
wire R7C16_GT00;
wire R3C45_GB00;
wire R20C33_GBO0;
wire R2C23_SPINE13;
wire R15C32_GB30;
wire R14C36_GB30;
wire R27C4_GB40;
wire R9C10_GB00;
wire R18C39_GB40;
wire R10C19_E20;
wire R5C25_GB20;
wire R1C1_A4;
wire R10C26_S83;
wire R6C22_GB30;
wire R28C25_CLK2;
wire R13C16_GB30;
wire R11C22_GB60;
wire R16C6_GT10;
wire R9C32_GB60;
wire R10C16_W21;
wire R7C15_GT00;
wire R16C35_GBO0;
wire R20C26_GT10;
wire R12C45_GB40;
wire R14C15_GB10;
wire R23C15_GB20;
wire R2C11_GBO0;
wire R22C42_GBO0;
wire R11C33_GB50;
wire R22C19_GT00;
wire R28C13_S26;
wire R3C31_GB20;
wire R18C15_GB00;
wire R24C9_GB70;
wire R1C28_W13;
wire R5C16_GB40;
wire R21C21_GBO0;
wire R10C19_SEL5;
wire R28C22_S80;
wire R23C20_GB60;
wire R7C45_GB00;
wire R12C27_GB30;
wire R12C2_GB40;
wire R25C35_GB00;
wire R10C37_B1;
wire R26C3_GB60;
wire R28C22_C1;
wire R20C14_GB00;
wire R28C31_Q2;
wire R26C7_GT00;
wire R22C46_GT10;
wire R25C4_GB20;
wire R27C12_GB00;
wire R22C25_GB40;
wire R2C20_GB30;
wire R23C31_GB20;
wire R26C22_GB70;
wire R11C21_GBO0;
wire R25C9_GT10;
wire R18C36_GBO1;
wire R3C28_GB20;
wire R22C38_GB50;
wire R12C31_GB70;
wire R3C9_GB60;
wire R23C12_GB20;
wire R16C18_GT10;
wire R9C14_GB30;
wire R21C45_GB60;
wire R26C10_GBO0;
wire R15C38_GB70;
wire R11C18_GB40;
wire R28C7_F2;
wire R3C37_GB10;
wire R28C28_W24;
wire R16C36_GB30;
wire R23C41_GB00;
wire R10C27_S10;
wire R6C26_GBO0;
wire R13C26_GB40;
wire R4C13_GB30;
wire R11C43_GB70;
wire R21C5_GBO0;
wire R17C27_GB70;
wire R16C23_GB60;
wire R4C40_GBO1;
wire R16C38_GB50;
wire R28C4_B0;
wire R23C4_GT00;
wire R12C29_GB50;
wire R10C26_W81;
wire R15C37_GB50;
wire R4C27_GB00;
wire R29C28_S21;
wire R7C27_GB30;
wire R10C34_N81;
wire R18C15_GB20;
wire R10C19_E82;
wire R20C29_GT00;
wire R27C9_GB50;
wire R10C30_B5;
wire R8C5_GB20;
wire R8C22_GT00;
wire R8C35_GBO1;
wire R1C47_D1;
wire R13C3_GBO1;
wire R1C47_CLK2;
wire R10C25_CLK0;
wire R29C28_S25;
wire R11C4_GB60;
wire R7C8_GB20;
wire R4C7_GB00;
wire R10C28_W11;
wire R17C39_GT00;
wire R8C17_GB60;
wire R22C3_GBO1;
wire R10C10_F2;
wire R25C11_GB60;
wire R3C12_GB70;
wire R5C37_GT00;
wire R21C26_GB40;
wire R6C3_GB10;
wire R9C44_GB60;
wire R14C13_GB70;
wire R4C40_GB60;
wire R10C10_A4;
wire R10C43_C6;
wire R20C10_GBO0;
wire R10C25_E22;
wire R13C26_GB10;
wire R23C29_GBO0;
wire R3C42_GB50;
wire R10C19_D0;
wire R6C26_GB40;
wire R12C24_GB40;
wire R23C34_GB50;
wire R10C43_F6;
wire R21C21_GBO1;
wire R10C30_UNK127;
wire R14C40_GB50;
wire R28C10_CE0;
wire R8C22_GBO1;
wire R28C43_C3;
wire R10C10_F7;
wire R2C43_GT00;
wire R15C11_GT10;
wire R8C24_GT00;
wire R11C14_GBO0;
wire R27C3_GB50;
wire R8C41_GB50;
wire R4C42_GT10;
wire R27C29_GB60;
wire R10C31_S81;
wire R28C13_F3;
wire R9C46_GT10;
wire R16C16_GT00;
wire R14C40_GB40;
wire R14C22_GB30;
wire R8C3_GB30;
wire R23C12_GBO0;
wire R10C25_N21;
wire R28C19_EW10;
wire R14C7_GT00;
wire R10C22_D3;
wire R23C17_GT00;
wire R27C12_GB60;
wire R2C44_GB20;
wire R21C19_GB10;
wire R17C14_GB40;
wire R14C32_GB30;
wire R23C45_GT10;
wire R27C36_GB40;
wire R7C20_GT10;
wire R20C42_GB40;
wire R23C33_GBO1;
wire R12C33_GB50;
wire R20C38_GB70;
wire R24C26_GBO1;
wire R21C3_GB20;
wire R5C7_GB20;
wire R20C29_GBO1;
wire R10C28_N23;
wire R8C27_GT00;
wire R25C5_GB70;
wire R23C36_GB00;
wire R28C4_F3;
wire R22C24_GB10;
wire R28C25_E83;
wire R6C32_GT00;
wire R2C43_SPINE1;
wire R10C28_B3;
wire R21C46_GT00;
wire R18C25_GB70;
wire R9C4_GB60;
wire R27C43_GBO0;
wire R4C44_GB20;
wire R1C1_F4;
wire R28C37_A4;
wire R28C16_B6;
wire R3C45_GT10;
wire R11C2_GB50;
wire R9C9_GBO0;
wire R11C16_GT00;
wire R9C32_GB30;
wire R1C32_D0;
wire R28C46_E26;
wire R4C25_GB30;
wire R23C20_GBO1;
wire R28C43_N80;
wire R8C43_GB00;
wire R28C31_D0;
wire R9C29_GB10;
wire R14C22_GT00;
wire R6C45_GB60;
wire R28C28_N83;
wire R9C38_GBO0;
wire R15C19_GT00;
wire R17C30_GB50;
wire R7C15_GB00;
wire R10C28_W83;
wire R2C14_GT00;
wire R17C25_GB60;
wire R28C46_D2;
wire R8C34_GB00;
wire R17C14_GB10;
wire R18C30_GB50;
wire R28C16_D0;
wire R5C7_GT00;
wire R22C43_GT00;
wire R21C35_GB10;
wire R10C43_S11;
wire R18C33_GB40;
wire R12C46_GB40;
wire R9C8_GB10;
wire R18C40_GB40;
wire R1C47_X02;
wire R10C28_W13;
wire R10C31_X06;
wire R9C8_GB60;
wire R17C24_GT00;
wire R24C42_GB70;
wire R12C40_GB50;
wire R13C9_GBO0;
wire R18C46_GB40;
wire R8C38_GBO0;
wire R10C22_F4;
wire R10C30_S23;
wire R7C6_GT00;
wire R4C2_GBO0;
wire R13C22_GB10;
wire R3C9_GB30;
wire R27C44_GB30;
wire R1C47_S81;
wire R10C34_W27;
wire R22C42_GT00;
wire R3C6_GB00;
wire R10C34_N20;
wire R22C7_GB60;
wire R15C36_GBO0;
wire R9C29_GB50;
wire R28C4_B5;
wire R10C25_S82;
wire R10C25_X03;
wire R6C22_GBO0;
wire R16C22_GB50;
wire R23C10_GB40;
wire R21C9_GB70;
wire R8C43_GB60;
wire R28C16_E23;
wire R16C40_GB30;
wire R21C2_GB20;
wire R1C28_E13;
wire R7C35_GB00;
wire R10C28_N13;
wire R13C31_GB40;
wire R22C12_GBO0;
wire R14C35_GB60;
wire R25C5_GB40;
wire R3C34_GT00;
wire R21C24_GT00;
wire R26C1_GBO0;
wire R10C25_N26;
wire R17C13_GT10;
wire R23C46_GB10;
wire R18C8_GB20;
wire R20C4_SPINE20;
wire R26C25_GT00;
wire R14C39_GT00;
wire R28C25_D6;
wire R14C44_GB50;
wire R10C27_EW10;
wire R15C18_GB70;
wire R3C34_GB40;
wire R13C6_GB20;
wire R25C31_GB60;
wire R25C32_GB60;
wire R11C16_GB50;
wire R26C4_GT10;
wire R18C33_GBO1;
wire R18C42_GBO1;
wire R7C30_GBO1;
wire R6C35_GB70;
wire R2C18_GBO0;
wire R10C34_S21;
wire R6C32_GB60;
wire R10C27_B5;
wire R22C42_GT10;
wire R28C7_E22;
wire R25C21_GBO0;
wire R23C9_GB30;
wire R10C27_EW20;
wire R12C3_GB40;
wire R27C32_GB60;
wire R12C13_GT00;
wire R15C2_GBO1;
wire R26C1_GT10;
wire R6C21_GT00;
wire R24C12_GBO0;
wire R25C44_GB60;
wire R10C37_C0;
wire R9C4_GT00;
wire R15C12_GT00;
wire R16C35_GB70;
wire R7C41_GB10;
wire R11C46_GB60;
wire R23C5_GB10;
wire R21C20_GB60;
wire R28C43_SEL6;
wire R14C11_GB70;
wire R1C1_S20;
wire R2C13_GB40;
wire R10C25_W26;
wire R14C46_GT10;
wire R10C37_S27;
wire R27C21_GB10;
wire R24C22_GB60;
wire R24C26_GB60;
wire R23C15_GBO1;
wire R2C21_GB40;
wire R14C32_GB00;
wire R10C28_F1;
wire R22C43_GB50;
wire R28C4_E11;
wire R27C2_GBO0;
wire R25C33_GB50;
wire R10C22_D1;
wire R28C37_A6;
wire R5C39_GT10;
wire R17C32_GB00;
wire R12C17_GB50;
wire R15C17_GT00;
wire R4C8_GT00;
wire R7C12_GB70;
wire R14C15_GB20;
wire R17C35_GB10;
wire R13C1_GT00;
wire R29C28_E11;
wire R10C34_W80;
wire R1C1_E20;
wire R28C10_D4;
wire R7C27_GB10;
wire R10C22_N22;
wire R9C44_GB00;
wire R11C23_GB20;
wire R5C23_GB50;
wire R22C17_GBO0;
wire R4C28_GB10;
wire R24C12_GB70;
wire R10C16_W26;
wire R13C11_GB60;
wire R1C32_E80;
wire R12C11_GB20;
wire R6C24_GB00;
wire R3C39_GB10;
wire R4C11_GB40;
wire R12C22_GB20;
wire R24C8_GB50;
wire R23C30_GBO0;
wire R28C7_F3;
wire R28C16_W81;
wire R25C33_GB40;
wire R26C31_GT00;
wire R6C30_GB00;
wire R22C42_GB50;
wire R15C27_GB10;
wire R10C28_E24;
wire R18C13_GT10;
wire R18C39_GB70;
wire R10C27_SEL7;
wire R1C28_Q1;
wire R10C37_A5;
wire R1C32_X06;
wire R5C39_GB70;
wire R10C40_S13;
wire R21C41_GB60;
wire R10C16_W23;
wire R17C19_GT00;
wire R5C9_GBO0;
wire R3C26_GBO1;
wire R10C22_S25;
wire R26C22_GB60;
wire R9C13_GB20;
wire R27C5_GT00;
wire R10C37_Q7;
wire R28C43_E12;
wire R28C10_S23;
wire R21C41_GB20;
wire R13C7_GB10;
wire R2C22_GB00;
wire R22C25_GT00;
wire R2C3_GB20;
wire R1C32_E13;
wire R26C21_GT00;
wire R25C28_GB30;
wire R20C13_GB50;
wire R5C35_GB30;
wire R17C44_GB00;
wire R16C39_GBO0;
wire R17C37_GB70;
wire R28C22_E24;
wire R28C31_B0;
wire R23C46_GBO1;
wire R18C33_GB60;
wire R25C10_GB00;
wire R15C14_GB00;
wire R4C28_GB70;
wire R8C25_GBO0;
wire R28C16_S24;
wire R1C47_F1;
wire R28C46_S25;
wire R23C46_GT10;
wire R25C15_GB40;
wire R16C14_GB00;
wire R22C29_GB40;
wire R17C32_GT00;
wire R26C5_GB00;
wire R6C3_GB40;
wire R8C38_GB20;
wire R28C34_D0;
wire R3C27_GB30;
wire R10C7_F4;
wire R23C8_GB30;
wire R18C18_GB10;
wire R24C12_GB30;
wire R10C29_N22;
wire R10C40_S82;
wire R27C13_GB60;
wire R5C43_GB40;
wire R11C40_GBO0;
wire R10C43_B5;
wire R10C27_CLK0;
wire R12C44_GBO0;
wire R8C14_GB30;
wire R17C34_GBO1;
wire R9C17_GT00;
wire R10C37_E23;
wire R16C15_GBO1;
wire R25C19_GT10;
wire R9C41_GBO0;
wire R4C44_GBO1;
wire R23C11_GBO1;
wire R6C21_GB40;
wire R13C29_GT10;
wire R10C25_B7;
wire R23C11_GB00;
wire R27C32_GB20;
wire R1C28_B2;
wire R10C27_A6;
wire R28C10_E82;
wire R9C20_GB50;
wire R24C15_GT10;
wire R28C22_C3;
wire R3C21_GT00;
wire R2C14_GB20;
wire R22C18_GBO0;
wire R7C16_GB70;
wire R6C24_GT10;
wire R13C21_GB60;
wire R15C24_GB20;
wire R26C33_GBO0;
wire R10C34_Q7;
wire R2C20_SPINE8;
wire R15C4_GB30;
wire R12C12_GBO0;
wire R13C3_GT00;
wire R20C25_GB30;
wire R26C27_GB30;
wire R5C2_GT00;
wire R28C10_E21;
wire R18C45_GB20;
wire R13C14_GB70;
wire R10C19_X02;
wire R16C15_GB60;
wire R25C7_GT00;
wire R11C44_GT10;
wire R6C19_GB00;
wire R28C10_Q5;
wire R21C15_GB20;
wire R27C38_GB20;
wire R2C11_GB50;
wire R4C26_GT10;
wire R18C27_GB30;
wire R1C32_N80;
wire R28C37_E83;
wire R14C45_GT00;
wire R2C32_SPINE4;
wire R10C10_S26;
wire R15C46_GT00;
wire R4C8_GBO0;
wire R28C28_D4;
wire R24C25_GBO1;
wire R4C30_GB10;
wire R16C29_GB60;
wire R3C16_GB50;
wire R14C16_GB40;
wire R17C12_GT00;
wire R28C40_S21;
wire R16C43_GB50;
wire R1C1_Q0;
wire R2C23_GB70;
wire R13C40_GB60;
wire R27C15_GB00;
wire R20C4_GB00;
wire R28C37_A3;
wire R28C43_N81;
wire R14C24_GB40;
wire R3C7_GB50;
wire R5C24_GB10;
wire R14C33_GB50;
wire R14C19_GB10;
wire R24C14_GB30;
wire R18C18_GB60;
wire R15C21_GT00;
wire R1C1_EW10;
wire R10C40_S26;
wire R6C14_GB50;
wire R10C7_X03;
wire R10C26_SN10;
wire R25C34_GB00;
wire R2C31_GB00;
wire R16C46_GB10;
wire R23C41_GBO0;
wire R28C28_C1;
wire R8C8_GB70;
wire R23C30_GB50;
wire R24C8_GB00;
wire R12C25_GB00;
wire R6C5_GB50;
wire R28C43_N82;
wire R28C46_X07;
wire R25C10_GBO0;
wire R25C30_GB40;
wire R24C34_GB20;
wire R12C3_GB00;
wire R16C44_GB30;
wire R6C43_GB20;
wire R13C10_GT00;
wire R14C35_GB40;
wire R25C35_GB50;
wire R8C41_GB10;
wire R12C18_GB50;
wire R10C22_E24;
wire R28C40_B1;
wire R15C10_GBO1;
wire R16C36_GB00;
wire R10C28_N10;
wire R27C12_GB20;
wire R13C2_GB40;
wire R21C44_GT10;
wire R23C41_GT10;
wire R21C28_GB30;
wire R12C22_GB30;
wire R8C24_GB10;
wire R8C37_GB10;
wire R27C23_GT00;
wire R8C35_GT10;
wire R2C36_GB40;
wire R10C25_B2;
wire R4C30_GB60;
wire R11C34_GT00;
wire R14C8_GB10;
wire R11C12_GBO1;
wire R22C13_GT00;
wire R10C29_E10;
wire R12C30_GT00;
wire R8C3_GB20;
wire R2C40_GBO0;
wire R16C43_GB40;
wire R10C40_N20;
wire R8C34_GB20;
wire R16C31_GB10;
wire R2C39_GB20;
wire R4C23_GT00;
wire R6C33_GB60;
wire R26C26_GB20;
wire R12C30_GB60;
wire R14C32_GT10;
wire R9C18_GB00;
wire R6C26_GB00;
wire R1C32_E82;
wire R13C12_GBO1;
wire R22C2_GBO0;
wire R27C17_GB00;
wire R14C8_GB00;
wire R18C17_GB20;
wire R24C31_GB50;
wire R10C37_A6;
wire R28C4_Q0;
wire R28C4_N25;
wire R28C13_S80;
wire R29C28_W81;
wire R21C19_GT00;
wire R23C43_GB70;
wire R15C35_GBO1;
wire R7C30_GB70;
wire R5C31_GB30;
wire R24C23_GB30;
wire R23C2_GBO1;
wire R1C28_X06;
wire R17C13_GB10;
wire R10C27_Q2;
wire R29C28_S23;
wire R21C6_GB70;
wire R25C14_GB30;
wire R28C13_F0;
wire R21C35_GB60;
wire R7C29_GBO0;
wire R10C16_B0;
wire R13C45_GB30;
wire R15C45_GB60;
wire R16C12_GB10;
wire R11C33_GBO0;
wire R24C12_GBO1;
wire R10C22_B2;
wire R28C16_E20;
wire R15C35_GB70;
wire R26C29_GB60;
wire R18C21_GB10;
wire R12C36_GB60;
wire R10C30_F1;
wire R15C30_GBO1;
wire R10C10_B6;
wire R10C37_E25;
wire R28C7_CE0;
wire R21C17_GT00;
wire R5C42_GB30;
wire R6C9_GB10;
wire R3C10_GBO0;
wire R23C13_GB30;
wire R6C4_GT10;
wire R2C28_GB70;
wire R12C10_GB30;
wire R7C10_GB50;
wire R15C24_GB50;
wire R20C35_GB10;
wire R16C38_GB70;
wire R10C22_X08;
wire R10C31_E81;
wire R10C29_SPINE26;
wire R21C22_GB10;
wire R24C8_GBO1;
wire R28C19_S11;
wire R21C11_GBO0;
wire R9C46_GB10;
wire R24C5_GB30;
wire R2C23_GT10;
wire R10C34_F4;
wire R10C34_N25;
wire R12C32_GB00;
wire R7C5_GB10;
wire R9C19_GB00;
wire R2C40_GB10;
wire R28C4_E24;
wire R2C5_GB20;
wire R1C32_D4;
wire R25C8_GB50;
wire R24C6_GB10;
wire R10C30_X08;
wire R10C30_F0;
wire R21C23_GBO0;
wire R3C32_GBO1;
wire R25C30_GB60;
wire R1C47_Q6;
wire R28C22_E20;
wire R9C13_GB60;
wire R6C31_GBO1;
wire R2C34_GB40;
wire R13C18_GB30;
wire R1C32_S12;
wire R21C39_GB00;
wire R6C27_GB30;
wire R22C9_GB60;
wire R28C7_N12;
wire R17C45_GB30;
wire R18C37_GT00;
wire R11C23_GBO0;
wire R8C46_GB00;
wire R17C43_GB50;
wire R10C16_N21;
wire R28C22_C4;
wire R16C11_GB10;
wire R15C32_GB60;
wire R9C29_GT10;
wire R20C46_GB70;
wire R11C8_GB20;
wire R1C32_LSR2;
wire R9C18_GB40;
wire R6C15_GB30;
wire R20C30_GB00;
wire R10C28_C7;
wire R1C28_C7;
wire R22C16_GB00;
wire R14C3_GB60;
wire R7C1_GT00;
wire R10C27_N26;
wire R8C12_GT00;
wire R1C1_D6;
wire R17C46_GB40;
wire R3C40_GB50;
wire R10C30_A1;
wire R28C46_C4;
wire R7C34_GT10;
wire R3C43_GT00;
wire R18C31_GT00;
wire R25C14_GB20;
wire R20C12_GB10;
wire R10C30_W22;
wire R3C31_GT00;
wire R15C3_GB70;
wire R9C45_GBO1;
wire R18C20_GB20;
wire R27C3_GBO1;
wire R8C32_GBO0;
wire R4C35_GB00;
wire R25C43_GB40;
wire R25C41_GB60;
wire R10C19_N22;
wire R28C19_LSR2;
wire R9C30_GB60;
wire R26C11_GB60;
wire R28C13_F5;
wire R28C10_W80;
wire R13C36_GB30;
wire R28C37_S22;
wire R28C4_A1;
wire R1C1_C4;
wire R22C46_GT00;
wire R5C35_GB20;
wire R24C13_GB40;
wire R22C15_GB60;
wire R1C32_CE1;
wire R28C19_S27;
wire R9C21_GT10;
wire R26C36_GT00;
wire R28C37_SEL0;
wire R25C27_GB70;
wire R22C41_GT00;
wire R13C30_GB50;
wire R28C34_S27;
wire R8C10_GB10;
wire R15C19_GB20;
wire R18C44_GBO0;
wire R13C25_GB70;
wire R10C7_W23;
wire R14C37_GBO1;
wire R6C13_GB00;
wire R10C29_SPINE25;
wire R3C17_GBO1;
wire R15C3_GB30;
wire R10C10_C7;
wire R21C10_GB70;
wire R2C44_GB00;
wire R6C37_GB20;
wire R18C7_GT10;
wire R25C20_GB40;
wire R9C32_GBO0;
wire R4C45_GB40;
wire R17C5_GB10;
wire R15C34_GB60;
wire R18C46_GB60;
wire R10C19_N12;
wire R20C25_GB70;
wire R3C35_GBO1;
wire R9C44_GB50;
wire R24C13_GB70;
wire R28C13_C6;
wire R15C25_GB10;
wire R28C19_W83;
wire R21C42_GB20;
wire R10C16_B2;
wire R28C31_C3;
wire R14C25_GT10;
wire R28C19_SEL5;
wire R21C13_GB30;
wire R20C15_GB50;
wire R10C27_W83;
wire R22C44_GB20;
wire R3C33_GB20;
wire R10C22_D7;
wire R10C22_W21;
wire R28C31_A0;
wire R12C29_GBO1;
wire R10C25_N24;
wire R5C24_GB40;
wire R14C35_GB30;
wire R28C34_S25;
wire R28C37_LSR1;
wire R11C29_GB10;
wire R1C28_E27;
wire R28C25_A2;
wire R28C46_N23;
wire R7C2_GT10;
wire R22C4_GB60;
wire R21C32_GB10;
wire R21C7_GB10;
wire R4C5_GB70;
wire R8C35_GB40;
wire R1C47_X05;
wire R28C4_SEL0;
wire R24C44_GB10;
wire R7C46_GT00;
wire R28C10_E24;
wire R14C24_GB10;
wire R6C39_GT00;
wire R8C16_GBO1;
wire R24C17_GB60;
wire R3C37_GBO0;
wire R28C25_B1;
wire R28C19_A0;
wire R7C27_GB00;
wire R18C14_GB20;
wire R16C38_GB10;
wire R2C10_GBO1;
wire R25C45_GB00;
wire R28C7_S20;
wire R8C16_GB40;
wire R3C31_GBO0;
wire R29C28_B2;
wire R21C6_GB50;
wire R8C26_GB30;
wire R10C26_N82;
wire R29C28_W80;
wire R28C46_E24;
wire R21C22_GB60;
wire R5C21_GB70;
wire R21C7_GB70;
wire R13C11_GB10;
wire R18C20_GB00;
wire R7C44_GB70;
wire R9C13_GB50;
wire R2C24_GT10;
wire R14C10_GB30;
wire R28C40_Q4;
wire R11C12_GB00;
wire R8C16_GB20;
wire R25C13_GB00;
wire R17C21_GB50;
wire R2C36_GB70;
wire R10C28_N22;
wire R26C7_GB60;
wire R12C5_GB60;
wire R8C38_GT10;
wire R16C32_GB50;
wire R12C20_GB40;
wire R13C14_GBO1;
wire R13C2_GB60;
wire R28C34_W24;
wire R18C31_GT10;
wire R12C14_GB10;
wire R28C16_W22;
wire R28C19_E26;
wire R28C16_Q3;
wire R13C16_GT00;
wire R17C3_GB00;
wire R15C42_GB40;
wire R3C33_GB10;
wire R25C43_GB60;
wire R14C23_GB00;
wire R8C19_GB00;
wire R4C12_GT10;
wire R18C26_GB70;
wire R28C31_N27;
wire R22C14_GB50;
wire R8C35_GB50;
wire R7C26_GT10;
wire R23C11_GB40;
wire R14C5_GB60;
wire R5C44_GB70;
wire R20C16_GB60;
wire R27C33_GT00;
wire R4C23_GB70;
wire R14C11_GT10;
wire R14C3_GB30;
wire R15C21_GBO0;
wire R22C10_GB50;
wire R10C16_D3;
wire R12C15_GB40;
wire R8C35_GBO0;
wire R10C37_W82;
wire R23C23_GBO0;
wire R17C23_GT10;
wire R21C4_GB30;
wire R18C24_GB60;
wire R8C45_GB00;
wire R10C30_X07;
wire R7C4_GBO1;
wire R21C38_GB00;
wire R16C34_GBO1;
wire R12C44_GT00;
wire R28C7_W20;
wire R9C10_GBO1;
wire R3C9_GT00;
wire R17C11_GB30;
wire R28C13_N80;
wire R28C34_N12;
wire R2C28_GT00;
wire R3C26_GT00;
wire R2C17_GB40;
wire R6C27_GBO0;
wire R18C21_GB00;
wire R29C28_E22;
wire R24C18_GB10;
wire R9C10_GT10;
wire R23C13_GB40;
wire R7C31_GBO0;
wire R2C33_GB50;
wire R10C29_C0;
wire R8C36_GB70;
wire R17C42_GBO0;
wire R15C5_GB10;
wire R15C20_GB50;
wire R25C2_GB60;
wire R21C36_GB70;
wire R20C2_GT10;
wire R28C13_S83;
wire R1C1_B5;
wire R1C47_W83;
wire R10C43_W26;
wire R10C37_W25;
wire R23C40_GB20;
wire R25C8_GT10;
wire R8C16_GT10;
wire R6C32_GB00;
wire R26C40_GBO0;
wire R12C19_GB30;
wire R10C10_E24;
wire R10C30_A3;
wire R28C40_A1;
wire R28C37_F6;
wire R1C47_E81;
wire R25C13_GB40;
wire R10C29_N25;
wire R3C9_GT10;
wire R26C18_GT10;
wire R11C21_GB50;
wire R28C40_SN10;
wire R4C6_GB60;
wire R10C37_B4;
wire R16C6_GBO1;
wire R7C20_GB60;
wire R11C10_GBO0;
wire R29C28_W27;
wire R23C26_GT10;
wire R28C37_N24;
wire R7C3_GB00;
wire R3C6_GBO0;
wire R4C14_GB00;
wire R4C10_GBO0;
wire R23C1_GBO1;
wire R2C38_GB70;
wire R9C41_GBO1;
wire R13C23_GB30;
wire R4C13_GB60;
wire R28C40_Q6;
wire R16C15_GB30;
wire R2C14_GB30;
wire R22C17_GB70;
wire R10C25_B4;
wire R28C19_N11;
wire R8C9_GB40;
wire R24C13_GB00;
wire R27C9_GB10;
wire R28C10_A1;
wire R28C37_W83;
wire R21C4_GB20;
wire R7C30_GB60;
wire R10C22_N25;
wire R15C12_GBO0;
wire R28C19_Q1;
wire R17C2_GB60;
wire R4C9_GB10;
wire R15C29_GB40;
wire R29C28_W23;
wire R2C3_SPINE13;
wire R21C19_GB50;
wire R2C11_GB20;
wire R16C36_GT10;
wire R11C11_GB70;
wire R6C36_GB70;
wire R24C2_GBO0;
wire R10C16_SN20;
wire R28C25_N25;
wire R1C1_E13;
wire R21C16_GB00;
wire R9C16_GB30;
wire R18C42_GB20;
wire R25C11_GB10;
wire R25C35_GB40;
wire R23C38_GB30;
wire R3C40_GBO0;
wire R13C42_GB50;
wire R14C18_GB00;
wire R3C31_GB40;
wire R20C31_GB10;
wire R8C35_GT00;
wire R13C43_GB40;
wire R10C30_S24;
wire R10C43_E80;
wire R10C43_B2;
wire R28C25_E27;
wire R28C31_SEL1;
wire R28C31_N80;
wire R27C33_GB40;
wire R28C13_A7;
wire R28C31_EW10;
wire R10C37_S20;
wire R3C26_GB30;
wire R27C12_GBO0;
wire R10C19_B1;
wire R1C47_W82;
wire R26C4_GB20;
wire R10C27_A7;
wire R26C6_GB40;
wire R28C40_N81;
wire R25C17_GB00;
wire R22C22_GT00;
wire R16C21_GB50;
wire R14C6_GB50;
wire R20C32_GB10;
wire R26C10_GB10;
wire R9C17_GB70;
wire R15C8_GB50;
wire R28C46_N22;
wire R1C47_S11;
wire R5C17_GB70;
wire R23C30_GT00;
wire R10C22_SEL0;
wire R28C28_LSR2;
wire R26C21_GBO1;
wire R10C26_S27;
wire R23C37_GB70;
wire R10C31_X03;
wire R9C46_GB50;
wire R28C13_X05;
wire R7C46_GB60;
wire R12C45_GB00;
wire R10C7_S81;
wire R28C34_SEL4;
wire R14C42_GT10;
wire R12C6_GB10;
wire R17C33_GB40;
wire R23C42_GB30;
wire R23C21_GT10;
wire R24C16_GB50;
wire R20C11_GB70;
wire R27C13_GBO1;
wire R10C22_A6;
wire R28C43_W25;
wire R17C2_GBO0;
wire R4C2_GB70;
wire R13C40_GB00;
wire R10C31_E25;
wire R9C19_GB50;
wire R11C43_GB60;
wire R9C22_GB00;
wire R9C21_GT00;
wire R4C13_GB20;
wire R23C20_GT10;
wire R22C18_GB40;
wire R25C11_GBO1;
wire R10C29_F3;
wire R9C30_GB50;
wire R26C12_GB10;
wire R8C43_GBO1;
wire R21C21_GB30;
wire R4C37_GB70;
wire R10C37_X06;
wire R28C4_A7;
wire R28C34_W23;
wire R7C22_GB20;
wire R12C3_GT10;
wire R10C10_S10;
wire R10C40_F1;
wire R26C33_GB60;
wire R14C7_GB60;
wire R20C42_GB30;
wire R6C14_GBO1;
wire R27C20_GT10;
wire R17C4_GB20;
wire R14C36_GB70;
wire R24C37_GB10;
wire R12C15_GBO0;
wire R24C35_GT10;
wire R10C29_D4;
wire R22C39_GBO0;
wire R10C29_SEL6;
wire R11C26_GB30;
wire R24C27_GB60;
wire R6C39_GB50;
wire R2C43_GBO1;
wire R25C34_GB30;
wire R28C7_W80;
wire R28C28_D0;
wire R18C10_GB40;
wire R26C31_GBO1;
wire R12C2_GB30;
wire R28C4_N27;
wire R18C25_GB10;
wire R28C16_F0;
wire R23C2_GB60;
wire R5C42_GT10;
wire R7C23_GB00;
wire R22C5_GB40;
wire R14C32_GB50;
wire R10C7_SEL7;
wire R18C7_GB20;
wire R28C16_S10;
wire R20C44_GB70;
wire R13C15_GB20;
wire R7C44_GB60;
wire R17C10_GBO1;
wire R22C38_GB60;
wire R10C25_CE0;
wire R4C46_GB60;
wire R8C27_GBO0;
wire R12C2_GB10;
wire R26C9_GB60;
wire R10C30_N22;
wire R18C22_GBO1;
wire R13C44_GB40;
wire R3C7_GB70;
wire R16C42_GB50;
wire R18C42_GT10;
wire R1C1_LSR1;
wire R27C10_GB70;
wire R10C16_N81;
wire R10C31_LSR2;
wire R28C46_LSR0;
wire R5C29_GB70;
wire R8C14_GT10;
wire R27C42_GBO0;
wire R16C38_GT00;
wire R26C27_GB70;
wire R22C9_GBO1;
wire R8C3_GT00;
wire R22C41_GB10;
wire R26C21_GB30;
wire R10C27_E20;
wire R24C3_GB50;
wire R10C37_W80;
wire R14C26_GBO1;
wire R5C22_GB20;
wire R9C45_GB40;
wire R3C11_GB50;
wire R10C43_C3;
wire R6C14_GT00;
wire R13C17_GB40;
wire R18C19_GB30;
wire R26C36_GBO1;
wire R26C29_GBO1;
wire R7C26_GB30;
wire R9C33_GB60;
wire R25C25_GB60;
wire R6C39_GB30;
wire R10C16_X02;
wire R28C19_X07;
wire R11C4_GB70;
wire R15C46_GB70;
wire R7C18_GB20;
wire R21C26_GBO1;
wire R6C29_GB20;
wire R29C28_A7;
wire R17C21_GB20;
wire R20C9_GB20;
wire R22C23_GB30;
wire R6C33_GBO1;
wire R10C34_SEL6;
wire R6C10_GB20;
wire R21C8_GB10;
wire R28C34_E21;
wire R21C2_GBO1;
wire R18C10_GB20;
wire R3C28_GB50;
wire R17C6_GT00;
wire R25C25_GBO0;
wire R15C19_GB00;
wire R25C22_GB60;
wire R28C37_D4;
wire R13C7_GB60;
wire R14C15_GB50;
wire R26C8_GB70;
wire R6C5_GB30;
wire R26C13_GB10;
wire R10C34_SN10;
wire R1C32_SN10;
wire R28C28_LSR1;
wire R10C43_W12;
wire R21C3_GB10;
wire R28C34_F4;
wire R29C28_Q0;
wire R6C26_GBO1;
wire R10C27_W21;
wire R28C31_E13;
wire R2C4_GB00;
wire R5C22_GB40;
wire R3C5_GB60;
wire R21C20_GBO0;
wire R3C13_GB50;
wire R21C16_GB30;
wire R23C7_GB50;
wire R24C32_GB60;
wire R5C18_GB50;
wire R10C10_S23;
wire R10C29_EW10;
wire R10C34_W23;
wire R28C10_S27;
wire R25C4_GB60;
wire R10C16_X08;
wire R2C36_GB60;
wire R24C23_GB60;
wire R26C45_GT00;
wire R7C41_GB70;
wire R10C16_D6;
wire R7C37_GB30;
wire R17C9_GB50;
wire R27C6_GB60;
wire R29C28_EW10;
wire R10C7_N83;
wire R6C44_GBO0;
wire R10C30_X02;
wire R22C43_GB40;
wire R21C13_GB10;
wire R22C25_GB20;
wire R22C4_GBO1;
wire R14C45_GB00;
wire R23C23_GB60;
wire R2C39_GT00;
wire R28C31_E20;
wire R12C2_GB70;
wire R26C20_GBO1;
wire R23C42_GT10;
wire R7C26_GB60;
wire R1C1_X08;
wire R28C22_LSR2;
wire R8C18_GT10;
wire R9C19_GB40;
wire R23C5_GB30;
wire R7C36_GBO0;
wire R28C4_X04;
wire R16C23_GBO1;
wire R10C37_C7;
wire R29C28_CLK1;
wire R24C35_GBO1;
wire R11C32_GT10;
wire R10C34_X03;
wire R2C11_GB10;
wire R15C10_GB50;
wire R22C32_GB10;
wire R10C43_CE0;
wire R8C20_GT00;
wire R6C15_GB40;
wire R23C26_GBO1;
wire R18C39_GBO1;
wire R10C25_CE1;
wire R10C10_X02;
wire R28C34_S21;
wire R12C39_GB10;
wire R16C24_GB10;
wire R25C23_GBO1;
wire R4C11_GB70;
wire R10C37_CE0;
wire R4C5_GB10;
wire R4C14_GBO0;
wire R22C5_GB10;
wire R18C12_GB20;
wire R24C28_GT10;
wire R11C37_GT10;
wire R12C14_GBO0;
wire R17C45_GB10;
wire R26C41_GB50;
wire R28C7_LSR0;
wire R1C1_X02;
wire R11C32_GB50;
wire R27C35_GBO1;
wire R7C31_GB10;
wire R15C6_GB70;
wire R7C26_GBO1;
wire R17C18_GBO0;
wire R22C25_GB70;
wire R1C47_N11;
wire R10C30_N25;
wire R1C28_S20;
wire R10C43_W27;
wire R28C37_N12;
wire R15C16_GT10;
wire R20C2_GBO0;
wire R2C44_GT10;
wire R13C21_GB70;
wire R10C34_W22;
wire R5C3_GBO1;
wire R28C40_E27;
wire R12C39_GT00;
wire R12C2_GBO1;
wire R23C28_GT10;
wire R28C22_Q6;
wire R21C39_GB30;
wire R10C26_X05;
wire R10C27_N27;
wire R16C30_GB60;
wire R26C29_GB30;
wire R15C46_GB10;
wire R28C4_F2;
wire R15C17_GB00;
wire R11C18_GBO1;
wire R12C46_GB60;
wire R10C26_SEL3;
wire R10C27_SEL3;
wire R25C31_GB40;
wire R5C24_GBO0;
wire R10C27_W27;
wire R26C27_GBO0;
wire R15C37_GT00;
wire R2C32_SPINE0;
wire R10C7_LSR2;
wire R28C4_S27;
wire R13C39_GB10;
wire R20C9_GT00;
wire R5C28_GB60;
wire R21C4_GB70;
wire R23C46_GB40;
wire R17C37_GT00;
wire R1C1_EW20;
wire R7C20_GB00;
wire R22C10_GB00;
wire R21C27_GB40;
wire R6C2_GT10;
wire R15C29_GBO0;
wire R17C27_GB00;
wire R5C27_GB70;
wire R8C28_GT00;
wire R17C7_GB60;
wire R24C25_GT00;
wire R21C23_GB20;
wire R25C46_GB10;
wire R10C43_E22;
wire R9C40_GB70;
wire R28C25_N12;
wire R10C19_S27;
wire R17C34_GB20;
wire R28C25_W22;
wire R28C34_E24;
wire R25C39_GB20;
wire R10C16_Q3;
wire R16C6_GB50;
wire R23C43_GB60;
wire R10C34_F5;
wire R28C16_N13;
wire R22C5_GBO0;
wire R25C43_GBO0;
wire R28C22_S22;
wire R6C7_GB50;
wire R8C39_GB00;
wire R4C21_GB70;
wire R3C21_GB40;
wire R5C12_GB60;
wire R26C45_GB00;
wire R2C12_GB20;
wire R18C30_GB60;
wire R10C31_SEL1;
wire R7C44_GB10;
wire R11C11_GB60;
wire R28C16_E11;
wire R1C28_D2;
wire R10C29_SN20;
wire R7C27_GB70;
wire R18C31_GBO1;
wire R14C9_GB00;
wire R16C31_GBO0;
wire R24C4_GB20;
wire R1C28_A0;
wire R10C22_LSR1;
wire R22C8_GBO1;
wire R10C29_S23;
wire R20C37_GB60;
wire R28C28_CE2;
wire R27C2_GB60;
wire R8C43_GB70;
wire R7C7_GBO0;
wire R9C6_GB40;
wire R5C43_GT00;
wire R17C13_GBO0;
wire R4C14_GB20;
wire R10C13_N83;
wire R9C6_GBO0;
wire R28C34_N13;
wire R28C22_S83;
wire R12C32_GT00;
wire R20C35_GB60;
wire R25C29_GB40;
wire R6C13_GB20;
wire R16C6_GB40;
wire R10C7_S83;
wire R10C10_N10;
wire R28C16_S27;
wire R28C37_W80;
wire R10C37_W23;
wire R9C28_GB00;
wire R25C28_GT10;
wire R10C29_W10;
wire R8C2_GB00;
wire R4C46_GBO1;
wire R22C40_GB70;
wire R10C40_N26;
wire R10C31_W81;
wire R9C18_GT00;
wire R13C2_GT10;
wire R21C24_GT10;
wire R1C1_S25;
wire R24C43_GB70;
wire R13C8_GT00;
wire R2C10_GB00;
wire R28C19_S25;
wire R17C18_GBO1;
wire R22C31_GB20;
wire R21C31_GB30;
wire R7C13_GT00;
wire R8C6_GB60;
wire R18C3_GB40;
wire R16C41_GB30;
wire R8C33_GBO0;
wire R8C4_GB10;
wire R14C26_GB10;
wire R1C47_C7;
wire R25C43_GB70;
wire R10C37_A0;
wire R28C13_S11;
wire R28C46_N26;
wire R27C29_GB30;
wire R10C10_W81;
wire R8C42_GB10;
wire R10C40_X02;
wire R10C13_SN10;
wire R9C21_GBO0;
wire R4C46_GB70;
wire R14C4_GB70;
wire R23C42_GBO1;
wire R24C44_GBO0;
wire R10C28_SEL7;
wire R16C5_GBO1;
wire R6C19_GB20;
wire R2C30_GBO1;
wire R27C33_GBO0;
wire R1C1_A5;
wire R10C27_X04;
wire R6C20_GB70;
wire R12C4_GB30;
wire R7C30_GB10;
wire R22C29_GBO0;
wire R18C9_GB40;
wire R17C27_GB40;
wire R16C15_GB00;
wire R28C28_E25;
wire R21C16_GBO1;
wire R14C2_GB60;
wire R17C42_GB00;
wire R23C39_GB70;
wire R1C32_A7;
wire R8C29_GB20;
wire R10C31_CLK0;
wire R1C47_A1;
wire R3C11_GB00;
wire R28C43_W11;
wire R11C23_GB50;
wire R28C34_Q7;
wire R16C22_GT00;
wire R25C44_GB00;
wire R9C24_GB10;
wire R18C36_GB00;
wire R10C37_Q1;
wire R22C17_GT00;
wire R3C5_GB00;
wire R10C22_X01;
wire R10C34_N80;
wire R10C40_N22;
wire R16C25_GB50;
wire R28C25_F1;
wire R21C31_GB40;
wire R21C17_GB00;
wire R28C31_E10;
wire R15C28_GB20;
wire R13C44_GBO0;
wire R25C35_GB20;
wire R27C36_GB20;
wire R26C26_GB00;
wire R21C41_GT10;
wire R27C10_GB40;
wire R25C32_GB20;
wire R10C37_N27;
wire R28C16_S80;
wire R12C13_GB70;
wire R28C16_B0;
wire R28C4_X01;
wire R7C8_GB70;
wire R9C33_GB10;
wire R20C28_GB40;
wire R24C33_GBO0;
wire R27C45_GBO1;
wire R10C22_W26;
wire R12C10_GT10;
wire R20C23_SPINE21;
wire R8C2_GB40;
wire R9C41_GB00;
wire R26C19_GBO0;
wire R21C24_GB70;
wire R22C34_GBO0;
wire R10C43_CLK2;
wire R5C46_GT00;
wire R12C27_GB60;
wire R14C22_GB60;
wire R12C19_GB60;
wire R16C19_GB60;
wire R6C38_GB00;
wire R4C23_GBO0;
wire R10C26_S20;
wire R28C13_Q7;
wire R20C24_GBO1;
wire R29C28_N81;
wire R4C23_GT10;
wire R12C6_GB40;
wire R24C15_GBO1;
wire R28C31_E82;
wire R10C7_S10;
wire R25C20_GBO1;
wire R28C31_E81;
wire R10C22_A2;
wire R11C39_GB50;
wire R22C21_GB50;
wire R10C30_W83;
wire R2C41_GBO0;
wire R10C26_E82;
wire R2C26_GT10;
wire R18C15_GB60;
wire R8C14_GBO1;
wire R17C44_GB20;
wire R25C15_GBO0;
wire R4C37_GB50;
wire R13C8_GB40;
wire R26C25_GB40;
wire R1C1_C0;
wire R2C26_GB60;
wire R12C3_GB30;
wire R18C20_GT10;
wire R4C19_GT00;
wire R27C15_GBO1;
wire R27C17_GB40;
wire R7C13_GBO1;
wire R17C26_GT10;
wire R23C46_GB20;
wire R22C2_GB30;
wire R9C11_GB20;
wire R1C28_N13;
wire R27C7_GT00;
wire R16C30_GB50;
wire R10C29_E12;
wire R9C33_GBO0;
wire R28C46_A0;
wire R17C8_GB50;
wire R13C27_GB60;
wire R23C4_GB50;
wire R2C17_SPINE11;
wire R12C26_GB50;
wire R21C18_GBO0;
wire R5C26_GB00;
wire R28C10_W24;
wire R25C12_GBO0;
wire R8C29_GBO1;
wire R28C31_X02;
wire R12C2_GB20;
wire R26C25_GBO0;
wire R10C13_W27;
wire R5C18_GB70;
wire R28C22_E10;
wire R4C3_GT10;
wire R5C19_GBO0;
wire R6C7_GB70;
wire R14C1_GBO0;
wire R21C21_GB40;
wire R26C3_GBO1;
wire R17C43_GB00;
wire R7C6_GB60;
wire R23C12_GB60;
wire R2C38_GBO1;
wire R26C35_GBO0;
wire R25C10_GT00;
wire R26C41_GB30;
wire R15C35_GB60;
wire R22C44_GT00;
wire R9C18_GBO0;
wire R13C32_GB70;
wire R10C43_W22;
wire R6C9_GBO1;
wire R17C3_GB60;
wire R26C44_GB40;
wire R10C16_N20;
wire R10C37_C5;
wire R11C20_GT10;
wire R9C20_GB40;
wire R2C39_GT10;
wire R26C6_GB20;
wire R22C9_GB40;
wire R9C30_GB40;
wire R1C1_Q7;
wire R29C28_W82;
wire R7C43_GB50;
wire R18C19_GB40;
wire R27C36_GB50;
wire R27C13_GB40;
wire R17C16_GB50;
wire R28C7_CLK2;
wire R12C42_GBO1;
wire R28C4_E27;
wire R8C25_GBO1;
wire R11C17_GBO0;
wire R23C11_GB60;
wire R2C23_GBO1;
wire R15C9_GB20;
wire R10C25_C0;
wire R10C29_S12;
wire R2C27_GBO0;
wire R17C7_GT00;
wire R21C16_GB10;
wire R9C3_GB10;
wire R11C7_GB40;
wire R20C46_GB30;
wire R24C14_GB00;
wire R5C33_GB30;
wire R10C30_S12;
wire R3C27_GB20;
wire R20C27_GB00;
wire R24C19_GBO0;
wire R12C10_GB00;
wire R4C5_GB30;
wire R13C30_GB60;
wire R10C40_CE0;
wire R24C33_GB40;
wire R27C44_GBO0;
wire R2C44_GT00;
wire R10C16_E21;
wire R28C43_EW20;
wire R10C7_C5;
wire R21C23_GT10;
wire R10C30_E24;
wire R10C40_F4;
wire R25C6_GB60;
wire R1C47_C6;
wire R3C23_GB30;
wire R2C39_GB60;
wire R16C26_GB60;
wire R26C14_GT00;
wire R23C10_GBO0;
wire R10C13_Q0;
wire R8C42_GB70;
wire R10C16_W13;
wire R28C4_E22;
wire R22C33_GB60;
wire R9C44_GB30;
wire R10C30_W82;
wire R28C43_D3;
wire R12C15_GB30;
wire R28C31_W25;
wire R10C43_N83;
wire R9C25_GB10;
wire R28C7_F0;
wire R8C33_GB40;
wire R4C37_GT10;
wire R8C20_GB20;
wire R16C2_GT00;
wire R4C17_GB30;
wire R13C26_GBO0;
wire R26C21_GB60;
wire R22C22_GB00;
wire R3C22_GT10;
wire R24C27_GT10;
wire R10C26_SEL1;
wire R11C36_GB20;
wire R17C33_GT10;
wire R28C16_W82;
wire R4C5_GT10;
wire R3C34_GT10;
wire R25C1_GBO1;
wire R11C44_GBO0;
wire R1C28_S81;
wire R4C8_GB30;
wire R15C27_GB40;
wire R17C6_GBO1;
wire R13C45_GT00;
wire R11C33_GB70;
wire R13C42_GB70;
wire R10C40_X03;
wire R10C7_EW20;
wire R1C1_W80;
wire R28C43_SEL4;
wire R10C26_F5;
wire R11C10_GB30;
wire R20C31_GT00;
wire R1C28_Q7;
wire R10C37_W20;
wire R20C20_GB50;
wire R28C40_A5;
wire R22C32_GT10;
wire R3C27_GB50;
wire R5C5_GB20;
wire R27C39_GB20;
wire R23C34_GB70;
wire R8C40_GT10;
wire R13C15_GBO0;
wire R1C1_W12;
wire R6C30_GB10;
wire R6C6_GBO0;
wire R28C37_F1;
wire R22C38_GB20;
wire R11C3_GB00;
wire R27C31_GB50;
wire R14C30_GBO1;
wire R6C20_GB00;
wire R18C22_GB70;
wire R10C26_LSR1;
wire R17C20_GB30;
wire R23C8_GB40;
wire R25C40_GB70;
wire R1C47_N20;
wire R25C22_GT00;
wire R10C30_D1;
wire R12C12_GB60;
wire R28C19_W25;
wire R28C19_B6;
wire R14C5_GT00;
wire R7C29_GB30;
wire R16C46_GB30;
wire R22C25_GBO0;
wire R23C12_GT10;
wire R1C32_F1;
wire R5C42_GB20;
wire R25C39_GT00;
wire R14C38_GBO1;
wire R23C11_GB30;
wire R15C26_GB20;
wire R11C31_GB40;
wire R22C13_GT10;
wire R4C11_GB10;
wire R3C18_GB40;
wire R2C43_GB20;
wire R4C30_GBO1;
wire R28C28_N80;
wire R17C36_GT10;
wire R4C12_GB50;
wire R15C33_GB20;
wire R14C38_GB30;
wire R17C16_GB60;
wire R28C37_SEL4;
wire R4C42_GT00;
wire R8C45_GB70;
wire R13C13_GB00;
wire R10C43_C4;
wire R21C41_GBO0;
wire R17C7_GB50;
wire R21C33_GT10;
wire R2C5_GB50;
wire R4C18_GB20;
wire R3C32_GB30;
wire R24C42_GB40;
wire R7C24_GBO1;
wire R22C33_GBO1;
wire R2C21_GB00;
wire R23C37_GT00;
wire R5C33_GBO0;
wire R4C36_GB50;
wire R14C30_GB40;
wire R12C9_GB10;
wire R27C16_GB20;
wire R3C19_GB40;
wire R20C38_GT10;
wire R25C43_GB20;
wire R13C22_GT00;
wire R27C22_GB30;
wire R1C1_W27;
wire R28C40_W27;
wire R22C18_GT10;
wire R24C43_GB40;
wire R24C36_GB60;
wire R18C29_GB70;
wire R6C33_GB40;
wire R10C26_E83;
wire R28C37_E81;
wire R5C40_GB40;
wire R20C17_GB50;
wire R17C2_GBO1;
wire R15C6_GB00;
wire R4C12_GB10;
wire R13C35_GB40;
wire R5C14_GB00;
wire R28C4_E83;
wire R28C40_D7;
wire R11C25_GB30;
wire R2C9_GB40;
wire R10C40_S24;
wire R10C30_E26;
wire R10C16_E10;
wire R24C7_GT00;
wire R9C16_GB00;
wire R4C44_GT10;
wire R21C37_GT00;
wire R16C5_GB20;
wire R11C7_GB20;
wire R28C37_LSR0;
wire R28C31_F4;
wire R10C26_D4;
wire R4C2_GB50;
wire R28C7_A5;
wire R10C26_F1;
wire R9C9_GB50;
wire R9C23_GT10;
wire R18C11_GB50;
wire R5C44_GBO1;
wire R16C8_GB10;
wire R7C29_GBO1;
wire R9C14_GB60;
wire R28C4_N10;
wire R23C23_GB30;
wire R14C31_GB40;
wire R5C6_GB70;
wire R18C30_GT10;
wire R16C11_GB40;
wire R11C9_GT10;
wire R6C38_GB60;
wire R10C27_C0;
wire R28C16_D7;
wire R3C17_GT00;
wire R28C22_A0;
wire R18C23_GB60;
wire R18C34_GBO1;
wire R12C18_GB70;
wire R27C18_GB10;
wire R18C32_GBO1;
wire R5C40_GBO1;
wire R9C4_GB40;
wire R27C40_GBO1;
wire R15C5_GT00;
wire R9C11_GBO0;
wire R25C12_GB50;
wire R12C28_GB70;
wire R28C31_A6;
wire R12C8_GB50;
wire R28C13_E25;
wire R8C23_GB30;
wire R21C30_GBO1;
wire R28C31_C7;
wire R9C21_GB30;
wire R28C46_SEL6;
wire R3C43_GB40;
wire R18C33_GT10;
wire R10C40_W81;
wire R7C10_GB40;
wire R28C25_X03;
wire R2C34_GB30;
wire R2C36_GT10;
wire R23C44_GBO1;
wire R10C7_SEL6;
wire R13C20_GBO1;
wire R25C39_GB00;
wire R11C22_GT10;
wire R13C29_GB70;
wire R17C21_GB00;
wire R9C21_GB50;
wire R1C47_E22;
wire R17C4_GT10;
wire R10C13_C1;
wire R24C34_GB50;
wire R1C47_B0;
wire R10C27_B7;
wire R28C10_C6;
wire R28C37_S81;
wire R15C25_GB00;
wire R9C34_GB60;
wire R21C20_GT10;
wire R8C42_GB60;
wire R10C10_X01;
wire R18C17_GB50;
wire R18C29_GB50;
wire R15C28_GB70;
wire R11C37_GBO1;
wire R1C28_Q2;
wire R5C18_GBO1;
wire R15C38_GB30;
wire R21C10_GB10;
wire R25C17_GT00;
wire R28C25_F7;
wire R22C11_GB00;
wire R21C4_GT10;
wire R22C46_GB40;
wire R10C22_A5;
wire R8C37_GB00;
wire R2C24_GB20;
wire R16C32_GB40;
wire R15C20_GB30;
wire R20C4_GB70;
wire R28C28_A0;
wire R20C12_GBO0;
wire R1C1_F0;
wire R1C32_S13;
wire R2C29_GT10;
wire R26C33_GB20;
wire R10C40_S22;
wire R6C1_GT10;
wire R10C29_A7;
wire R14C34_GBO1;
wire R2C11_GB00;
wire R24C16_GB00;
wire R15C13_GB10;
wire R17C16_GB40;
wire R16C33_GB50;
wire R10C19_F7;
wire R4C34_GT00;
wire R17C44_GBO1;
wire R12C41_GB60;
wire R25C30_GB50;
wire R12C37_GBO1;
wire R10C13_W10;
wire R10C29_Q6;
wire R6C4_GBO1;
wire R12C18_GBO1;
wire R21C31_GB00;
wire R13C28_GB20;
wire R5C7_GB70;
wire R17C9_GB60;
wire R12C34_GB50;
wire R5C11_GBO1;
wire R5C4_GB40;
wire R11C2_GT00;
wire R17C40_GB60;
wire R5C5_GB40;
wire R28C40_E20;
wire R22C22_GB20;
wire R16C38_GB40;
wire R5C26_GB50;
wire R25C7_GT10;
wire R18C39_GB50;
wire R10C22_W10;
wire R21C46_GB60;
wire R9C8_GB30;
wire R8C28_GB30;
wire R17C7_GB30;
wire R14C22_GBO0;
wire R7C18_GB60;
wire R21C10_GB40;
wire R20C38_GB00;
wire R9C46_GB00;
wire R10C19_B2;
wire R10C10_W82;
wire R10C30_A6;
wire R28C7_B2;
wire R18C36_GB60;
wire R11C8_GBO1;
wire R20C39_GBO1;
wire R2C12_GBO0;
wire R25C18_GBO0;
wire R6C7_GBO1;
wire R21C2_GB00;
wire R21C18_GB60;
wire R1C32_N27;
wire R15C29_GB30;
wire R10C13_B3;
wire R25C34_GT10;
wire R28C4_CLK0;
wire R16C20_GBO1;
wire R20C43_GBO1;
wire R10C19_W23;
wire R10C43_N20;
wire R18C18_GBO1;
wire R10C10_LSR0;
wire R26C20_GB00;
wire R8C9_GB30;
wire R28C40_CLK2;
wire R17C20_GB60;
wire R28C46_A4;
wire R6C21_GT10;
wire R23C28_GB50;
wire R3C2_GBO1;
wire R17C36_GB50;
wire R24C40_GB60;
wire R26C2_GB10;
wire R9C10_GBO0;
wire R10C19_E23;
wire R13C2_GT00;
wire R5C16_GB70;
wire R10C29_N20;
wire R2C30_GB70;
wire R10C25_S20;
wire R11C4_GB20;
wire R13C13_GB40;
wire R15C26_GB30;
wire R28C19_W10;
wire R3C27_GB00;
wire R28C28_W25;
wire R15C6_GB30;
wire R6C46_GT00;
wire R15C16_GB30;
wire R15C22_GB50;
wire R7C37_GB10;
wire R28C16_W83;
wire R14C44_GBO0;
wire R22C10_GT00;
wire R11C27_GBO1;
wire R21C35_GB30;
wire R22C37_GB30;
wire R10C22_S27;
wire R6C9_GB70;
wire R23C32_GB20;
wire R10C27_E82;
wire R28C40_X01;
wire R15C13_GBO0;
wire R16C9_GB60;
wire R9C42_GB30;
wire R11C42_GB70;
wire R22C31_GB60;
wire R1C1_Q6;
wire R10C26_CLK1;
wire R23C38_GB60;
wire R27C2_GB20;
wire R28C46_S21;
wire R15C15_GB10;
wire R10C10_D7;
wire R25C35_GB60;
wire R10C7_B1;
wire R5C36_GB60;
wire R28C22_E26;
wire R28C40_E10;
wire R27C19_GBO1;
wire R28C7_W25;
wire R1C1_C5;
wire R10C7_N82;
wire R4C33_GB20;
wire R12C45_GB30;
wire R5C41_GB20;
wire R28C40_W25;
wire R20C15_GT10;
wire R27C5_GB30;
wire R9C17_GBO0;
wire R17C20_GT10;
wire R7C17_GB30;
wire R17C3_GB10;
wire R5C11_GB30;
wire R10C29_W22;
wire R10C30_F2;
wire R10C34_D7;
wire R14C12_GB00;
wire R20C22_GBO0;
wire R23C25_GBO0;
wire R11C6_GB50;
wire R22C33_GB20;
wire R22C41_GB50;
wire R10C26_N24;
wire R6C17_GB20;
wire R22C44_GT10;
wire R21C25_GB00;
wire R11C45_GBO1;
wire R12C42_GB60;
wire R18C20_GB50;
wire R25C4_GB70;
wire R7C40_GB50;
wire R10C7_E82;
wire R27C25_GB30;
wire R17C2_GB20;
wire R17C30_GB00;
wire R10C26_W21;
wire R16C35_GB60;
wire R28C19_N23;
wire R28C28_N11;
wire R9C33_GB00;
wire R11C34_GB00;
wire R3C17_GB50;
wire R5C41_GBO1;
wire R17C17_GBO0;
wire R18C12_GB60;
wire R5C19_GB60;
wire R16C14_GB50;
wire R26C11_GB30;
wire R24C45_GB50;
wire R28C10_S22;
wire R23C16_GB70;
wire R28C10_F6;
wire R28C28_D3;
wire R27C31_GBO0;
wire R2C36_GBO0;
wire R12C19_GT10;
wire R8C17_GT00;
wire R5C21_GBO0;
wire R5C27_GB30;
wire R21C13_GB40;
wire R21C30_GB70;
wire R9C15_GB10;
wire R5C7_GBO1;
wire R20C33_GB00;
wire R10C28_S22;
wire R28C46_CLK2;
wire R10C34_B4;
wire R10C7_N22;
wire R5C45_GB40;
wire R1C1_CE1;
wire R22C21_GB40;
wire R15C35_GBO0;
wire R16C25_GB00;
wire R15C17_GB20;
wire R14C39_GT10;
wire R20C20_GB20;
wire R28C13_X02;
wire R16C10_GB50;
wire R10C19_E12;
wire R17C25_GB40;
wire R12C9_GBO1;
wire R25C4_GBO1;
wire R24C33_GT10;
wire R2C35_GB30;
wire R7C29_GB40;
wire R9C43_GBO1;
wire R22C35_GB10;
wire R25C9_GT00;
wire R15C33_GT00;
wire R1C47_S13;
wire R10C13_B2;
wire R16C28_GB70;
wire R28C31_S24;
wire R24C5_GB10;
wire R14C37_GB20;
wire R26C19_GB20;
wire R14C40_GB30;
wire R13C14_GB40;
wire R10C16_N24;
wire R11C15_GB00;
wire R22C31_GBO1;
wire R10C27_X07;
wire R28C16_D3;
wire R22C37_GB20;
wire R12C27_GB20;
wire R15C33_GB50;
wire R28C28_E27;
wire R18C33_GBO0;
wire R28C31_S21;
wire R2C13_GB50;
wire R7C29_GT10;
wire R9C37_GB60;
wire R14C38_GB00;
wire R4C30_GB30;
wire R11C16_GB40;
wire R13C39_GB30;
wire R13C43_GB60;
wire R22C15_GBO1;
wire R10C7_CLK2;
wire R10C16_S10;
wire R14C3_GB10;
wire R15C4_GBO0;
wire R6C20_GB60;
wire R27C40_GB60;
wire R9C2_GB40;
wire R8C41_GBO1;
wire R21C6_GBO0;
wire R3C24_GB60;
wire R10C13_N24;
wire R4C20_GT10;
wire R6C46_GB60;
wire R23C3_GT10;
wire R10C10_S13;
wire R28C10_E26;
wire R23C30_GBO1;
wire R25C10_GB20;
wire R28C4_LSR2;
wire R10C26_W26;
wire R18C14_GB10;
wire R24C16_GB10;
wire R28C43_LSR1;
wire R28C34_C3;
wire R23C33_GB10;
wire R13C36_GB10;
wire R1C32_B0;
wire R8C16_GT00;
wire R5C28_GB10;
wire R16C44_GT00;
wire R10C7_S21;
wire R12C26_GB40;
wire R25C22_GB10;
wire R16C8_GB00;
wire R13C18_GB40;
wire R13C6_GB50;
wire R28C4_D0;
wire R1C28_X05;
wire R1C1_SEL4;
wire R23C17_GBO0;
wire R7C41_GT00;
wire R9C42_GB10;
wire R6C20_GB30;
wire R15C16_GB50;
wire R10C31_W11;
wire R28C46_CLK0;
wire R28C43_S27;
wire R4C8_GB20;
wire R20C2_GB70;
wire R28C10_X03;
wire R1C32_W11;
wire R9C8_GT10;
wire R10C40_E20;
wire R20C43_GB00;
wire R28C13_W80;
wire R16C29_GBO0;
wire R27C39_GB00;
wire R20C40_GB60;
wire R22C34_GB70;
wire R28C43_S83;
wire R24C21_GB30;
wire R16C44_GB10;
wire R28C22_X06;
wire R10C29_UNK125;
wire R9C1_GT10;
wire R10C40_SEL1;
wire R28C16_X06;
wire R27C3_GB10;
wire R1C1_N82;
wire R21C46_GB50;
wire R15C30_GB30;
wire R15C40_GB60;
wire R9C5_GBO0;
wire R10C40_Q1;
wire R23C10_GT10;
wire R9C36_GB50;
wire R2C11_SPINE9;
wire R3C18_GB50;
wire R16C33_GB30;
wire R9C4_GB50;
wire R10C37_D5;
wire R21C7_GT10;
wire R25C24_GB50;
wire R12C33_GB60;
wire R24C19_GB30;
wire R10C34_W24;
wire R17C36_GB10;
wire R10C28_C0;
wire R11C35_GB50;
wire R28C4_LSR1;
wire R28C19_F1;
wire R2C16_GB50;
wire R26C8_GBO0;
wire R9C43_GB40;
wire R20C20_GB10;
wire R11C3_GB40;
wire R7C46_GB20;
wire R12C16_GBO0;
wire R28C22_SEL7;
wire R17C16_GB70;
wire R21C30_GB30;
wire R15C34_GBO1;
wire R23C8_GB10;
wire R26C38_GB30;
wire R11C23_GB00;
wire R21C8_GB40;
wire R9C6_GB00;
wire R10C27_N23;
wire R7C40_GT00;
wire R25C2_GB50;
wire R12C17_GB10;
wire R18C24_GT10;
wire R9C46_GT00;
wire R22C11_GB20;
wire R12C41_GB30;
wire R11C31_GB70;
wire R10C31_SEL2;
wire R12C7_GB30;
wire R5C20_GB40;
wire R10C19_CLK2;
wire R2C12_SPINE12;
wire R27C4_GB20;
wire R20C45_GB50;
wire R7C28_GB50;
wire R20C25_GB00;
wire R8C27_GB50;
wire R10C13_F2;
wire R7C6_GB30;
wire R27C5_GB70;
wire R21C39_GBO1;
wire R15C11_GB60;
wire R13C17_GB50;
wire R22C36_GB00;
wire R27C12_GB10;
wire R20C9_GB60;
wire R26C45_GBO1;
wire R6C16_GB00;
wire R20C45_GBO0;
wire R10C34_S26;
wire R20C23_GB10;
wire R4C33_GB50;
wire R11C33_GBO1;
wire R10C37_S22;
wire R12C25_GB20;
wire R2C18_GT10;
wire R23C45_GB50;
wire R4C11_GBO1;
wire R8C36_GBO0;
wire R12C14_GB70;
wire R21C38_GB40;
wire R2C40_GBO1;
wire R16C25_GBO0;
wire R10C43_LSR2;
wire R6C9_GB20;
wire R28C7_F6;
wire R11C23_GBO1;
wire R26C35_GB60;
wire R2C39_GBO0;
wire R24C19_GT10;
wire R15C4_GB00;
wire R22C19_GB00;
wire R12C36_GB30;
wire R10C26_N25;
wire R22C28_GB10;
wire R28C40_B4;
wire R10C27_B1;
wire R28C22_Q4;
wire R7C24_GB30;
wire R12C37_GB50;
wire R2C27_GT00;
wire R2C31_GBO0;
wire R9C42_GB20;
wire R21C34_GBO1;
wire R27C36_GB70;
wire R10C37_CLK0;
wire R28C19_N26;
wire R25C5_GBO1;
wire R11C40_GB00;
wire R23C16_GT10;
wire R25C11_GT10;
wire R20C15_GB30;
wire R11C28_GB70;
wire R7C5_GT00;
wire R12C44_GB10;
wire R8C11_GB30;
wire R10C37_F1;
wire R9C47_F6;
wire R17C36_GB40;
wire R28C31_N23;
wire R18C13_GB30;
wire R10C13_S11;
wire R28C43_S82;
wire R25C19_GB00;
wire R25C43_GB00;
wire R2C9_GB30;
wire R11C46_GB40;
wire R8C24_GT10;
wire R20C12_SPINE16;
wire R15C1_F6;
wire R21C39_GBO0;
wire R15C30_GB40;
wire R4C35_GB40;
wire R21C44_GB40;
wire R14C11_GB20;
wire R20C29_GB70;
wire R25C31_GBO0;
wire R12C7_GBO1;
wire R25C42_GB50;
wire R10C34_F1;
wire R28C25_D7;
wire R14C7_GBO1;
wire R10C28_D2;
wire R28C40_B5;
wire R23C3_GB00;
wire R10C40_W83;
wire R13C3_GB00;
wire R27C28_GB30;
wire R10C43_B1;
wire R27C3_GB40;
wire R1C1_S80;
wire R18C41_GT00;
wire R24C6_GT00;
wire R8C17_GB30;
wire R13C22_GB20;
wire R22C32_GT00;
wire R1C47_X07;
wire R13C3_GBO0;
wire R10C13_N27;
wire R28C19_X06;
wire R14C8_GB30;
wire R28C28_N26;
wire R5C14_GB10;
wire R12C42_GT10;
wire R14C35_GB50;
wire R28C4_E80;
wire R3C39_GT10;
wire R14C14_GB00;
wire R3C10_GB50;
wire R10C27_CE1;
wire R9C22_GT10;
wire R20C41_GBO0;
wire R4C32_GB70;
wire R26C14_GB00;
wire R24C28_GB20;
wire R10C7_Q1;
wire R28C4_S12;
wire R7C24_GB50;
wire R20C20_GB30;
wire R5C9_GB50;
wire R3C24_GB20;
wire R13C29_GB00;
wire R8C19_GB10;
wire R10C16_A3;
wire R21C24_GB00;
wire R24C2_GB10;
wire R23C22_GB70;
wire R14C17_GB60;
wire R12C33_GB00;
wire R1C1_C6;
wire R22C46_GB60;
wire R10C29_C5;
wire R11C35_GB30;
wire R10C30_SEL5;
wire R28C10_Q6;
wire R17C34_GB60;
wire R28C31_W23;
wire R26C18_GB00;
wire R11C12_GB50;
wire R17C5_GB20;
wire R23C17_GB10;
wire R26C8_GBO1;
wire R1C1_D7;
wire R29C28_CE0;
wire R13C44_GB60;
wire R28C46_D1;
wire R10C43_S27;
wire R26C9_GB10;
wire R10C26_D6;
wire R18C8_GB30;
wire R4C4_GT00;
wire R20C6_GB20;
wire R5C28_GB30;
wire R15C29_GT00;
wire R7C43_GBO0;
wire R14C34_GB70;
wire R20C15_GB00;
wire R10C27_CLK2;
wire R26C10_GT00;
wire R11C32_GBO0;
wire R17C13_GB00;
wire R15C17_GBO1;
wire R8C41_GB00;
wire R9C14_GB20;
wire R10C10_N20;
wire R27C24_GB10;
wire R1C47_Q3;
wire R10C30_C0;
wire R10C40_A0;
wire R12C37_GB60;
wire R13C30_GB10;
wire R5C4_GB20;
wire R23C20_GB10;
wire R25C7_GB30;
wire R8C39_GT10;
wire R17C23_GB50;
wire R15C35_GT10;
wire R16C45_GB10;
wire R10C10_B4;
wire R10C28_X06;
wire R28C34_E25;
wire R3C17_GB70;
wire R2C13_GBO0;
wire R5C27_GB50;
wire R14C18_GBO1;
wire R14C35_GBO0;
wire R26C18_GB50;
wire R26C4_GBO1;
wire R21C15_GBO0;
wire R22C4_GB40;
wire R27C32_GT10;
wire R1C47_W11;
wire R10C25_SEL3;
wire R21C4_GB10;
wire R14C34_GT00;
wire R10C43_W23;
wire R25C17_GB60;
wire R28C25_EW20;
wire R9C30_GT00;
wire R10C13_CE1;
wire R27C15_GB70;
wire R7C32_GB70;
wire R26C12_GT00;
wire R26C45_GB30;
wire R27C40_GB50;
wire R3C2_GB10;
wire R14C39_GB70;
wire R17C37_GBO0;
wire R26C19_GBO1;
wire R18C10_GB30;
wire R11C19_GB10;
wire R28C22_N22;
wire R28C34_W27;
wire R17C30_GB70;
wire R10C37_X01;
wire R27C20_GB60;
wire R26C31_GT10;
wire R4C45_GB20;
wire R7C16_GB20;
wire R1C1_SEL0;
wire R13C10_GB70;
wire R9C9_GB00;
wire R24C37_GT00;
wire R13C27_GB10;
wire R10C31_B0;
wire R21C27_GT00;
wire R2C27_GB10;
wire R13C27_GB20;
wire R10C7_E83;
wire R6C21_GB10;
wire R18C36_GT00;
wire R10C29_Q0;
wire R28C16_N12;
wire R26C24_GT10;
wire R1C32_EW20;
wire R4C43_GB60;
wire R7C44_GB40;
wire R9C29_GB20;
wire R2C43_SPINE5;
wire R7C34_GB40;
wire R23C21_GB10;
wire R16C9_GB70;
wire R23C41_GBO1;
wire R16C5_GB00;
wire R3C32_GB70;
wire R28C28_Q0;
wire R28C37_W81;
wire R13C46_GB30;
wire R3C20_GBO1;
wire R5C29_GB60;
wire R21C32_GB30;
wire R10C34_F0;
wire R28C4_F0;
wire R8C39_GBO0;
wire R8C3_GBO0;
wire R10C10_E83;
wire R27C23_GB10;
wire R24C38_GBO1;
wire R3C19_GBO1;
wire R22C18_GB50;
wire R10C16_B7;
wire R3C41_GB10;
wire R23C32_GB70;
wire R20C42_GBO0;
wire R5C7_GB60;
wire R7C43_GT00;
wire R24C2_GB20;
wire R17C26_GB20;
wire R16C13_GB50;
wire R25C38_GB30;
wire R10C13_CLK0;
wire R28C19_W21;
wire R13C9_GT10;
wire R10C29_N80;
wire R3C18_GBO0;
wire R14C14_GB60;
wire R17C18_GB40;
wire R16C30_GB00;
wire R15C34_GB20;
wire R13C18_GBO1;
wire R28C46_S22;
wire R23C21_GBO0;
wire R6C33_GB20;
wire R11C40_GB40;
wire R15C13_GB20;
wire R22C13_GB20;
wire R6C20_GB10;
wire R11C9_GB70;
wire R10C25_B3;
wire R16C5_GB60;
wire R11C30_GB50;
wire R10C25_A5;
wire R8C4_GBO1;
wire R7C21_GBO1;
wire R23C16_GB40;
wire R25C19_GBO0;
wire R8C28_GB00;
wire R8C43_GBO0;
wire R23C25_GB50;
wire R7C37_GT00;
wire R20C17_GB40;
wire R10C31_E24;
wire R8C44_GT00;
wire R24C20_GB30;
wire R10C37_S10;
wire R21C23_GB40;
wire R8C43_GB40;
wire R23C33_GB70;
wire R4C2_GB40;
wire R1C47_A5;
wire R10C7_Q0;
wire R28C19_C4;
wire R12C36_GB70;
wire R28C43_N83;
wire R12C8_GB20;
wire R17C13_GB40;
wire R14C19_GB30;
wire R9C39_GB00;
wire R25C40_GT10;
wire R9C3_GB00;
wire R2C39_GB40;
wire R15C30_GB60;
wire R28C40_C6;
wire R29C28_E10;
wire R27C25_GB20;
wire R15C42_GBO1;
wire R10C16_W82;
wire R10C27_Q0;
wire R16C29_GB70;
wire R2C6_GBO1;
wire R24C5_GBO0;
wire R16C17_GB60;
wire R6C36_GB60;
wire R26C35_GBO1;
wire R23C18_GBO0;
wire R15C20_GB70;
wire R18C6_GB50;
wire R23C36_GB50;
wire R2C29_GB60;
wire R10C34_D4;
wire R1C1_S22;
wire R8C6_GBO1;
wire R8C45_GBO1;
wire R10C13_A1;
wire R27C31_GB10;
wire R28C37_C4;
wire R16C11_GB00;
wire R15C4_GB20;
wire R9C23_GB10;
wire R12C20_GB50;
wire R23C24_GB10;
wire R3C18_GT10;
wire R21C11_GT00;
wire R11C31_GT10;
wire R11C20_GB20;
wire R15C43_GB20;
wire R24C43_GB30;
wire R16C28_GB50;
wire R10C19_W27;
wire R10C31_S27;
wire R10C40_W24;
wire R20C24_GB30;
wire R28C31_E23;
wire R14C1_GT00;
wire R1C1_B1;
wire R18C7_GB30;
wire R21C43_GBO1;
wire R2C10_GT00;
wire R29C28_S10;
wire R28C43_B5;
wire R28C28_E11;
wire R17C8_GT00;
wire R10C25_W10;
wire R1C47_N24;
wire R5C13_GB70;
wire R6C7_GB60;
wire R26C22_GB00;
wire R16C35_GB50;
wire R15C7_GBO1;
wire R12C19_GB40;
wire R5C44_GB00;
wire R7C33_GB20;
wire R28C4_SN20;
wire R11C10_GB20;
wire R14C23_GB30;
wire R27C28_GT00;
wire R1C1_SEL2;
wire R1C1_SEL3;
wire R10C25_S10;
wire R28C10_W83;
wire R10C30_SN20;
wire R20C29_GB10;
wire R17C35_GB20;
wire R11C25_GB20;
wire R1C47_X06;
wire R15C46_GB00;
wire R13C43_GB20;
wire R28C19_E82;
wire R10C28_UNK124;
wire R18C23_GT10;
wire R18C7_GB50;
wire R10C43_C0;
wire R28C34_N23;
wire R11C37_GB20;
wire R27C23_GB60;
wire R11C40_GB30;
wire R28C25_SEL7;
wire R28C16_Q2;
wire R8C21_GB10;
wire R28C13_F4;
wire R10C26_E22;
wire R10C30_C3;
wire R5C44_GT10;
wire R4C3_GB00;
wire R9C34_GT00;
wire R16C46_GB70;
wire R29C28_X05;
wire R2C39_GB70;
wire R13C13_GT10;
wire R16C19_GB10;
wire R12C18_GBO0;
wire R9C15_GB70;
wire R10C10_S12;
wire R15C11_GB20;
wire R20C45_GB70;
wire R29C28_N12;
wire R4C17_GB60;
wire R1C32_S20;
wire R28C10_X07;
wire R17C17_GB50;
wire R28C31_X04;
wire R2C11_GT10;
wire R2C30_GB20;
wire R10C7_Q6;
wire R12C23_GB20;
wire R6C22_GB50;
wire R28C46_EW20;
wire R22C28_GB00;
wire R10C29_C6;
wire R29C28_D4;
wire R10C7_C4;
wire R9C35_GBO0;
wire R11C36_GBO0;
wire R4C45_GB30;
wire R16C28_GB30;
wire R6C18_GB20;
wire R28C7_E27;
wire R27C9_GB00;
wire R7C33_GBO1;
wire R15C45_GB30;
wire R10C10_A7;
wire R10C25_X02;
wire R21C36_GBO0;
wire R9C31_GB20;
wire R20C25_GBO1;
wire R10C13_E22;
wire R10C29_W82;
wire R10C7_W81;
wire R9C31_GBO1;
wire R10C16_W25;
wire R10C27_N20;
wire R10C25_D4;
wire R28C7_W81;
wire R28C13_B5;
wire R4C16_GB40;
wire R28C13_W13;
wire R4C17_GT10;
wire R10C40_N21;
wire R27C2_GB00;
wire R4C28_GB60;
wire R17C33_GB70;
wire R7C3_GB70;
wire R10C29_SPINE29;
wire R3C19_GB20;
wire R4C31_GB70;
wire R1C32_N82;
wire R24C22_GT00;
wire R11C15_GB20;
wire R25C31_GB10;
wire R10C10_SEL2;
wire R16C30_GB70;
wire R8C30_GT10;
wire R10C27_E21;
wire R24C3_GBO0;
wire R11C9_GBO1;
wire R28C16_C3;
wire R9C13_GB70;
wire R10C10_Q5;
wire R28C13_LSR1;
wire R12C44_GB40;
wire R17C9_GB10;
wire R10C10_E81;
wire R10C34_N27;
wire R22C21_GT10;
wire R28C46_F5;
wire R2C27_GB50;
wire R15C36_GB70;
wire R10C16_LSR0;
wire R6C44_GBO1;
wire R18C19_GBO1;
wire R4C19_GB70;
wire R4C19_GT10;
wire R16C2_GB10;
wire R9C40_GBO1;
wire R17C2_GT00;
wire R21C39_GB20;
wire R17C24_GB00;
wire R22C7_GBO1;
wire R10C27_S20;
wire R10C31_D6;
wire R15C22_GT10;
wire R7C5_GB40;
wire R25C2_GBO1;
wire R7C40_GB60;
wire R14C43_GB10;
wire R26C25_GB00;
wire R2C28_GB40;
wire R12C24_GBO1;
wire R16C41_GB40;
wire R8C31_GBO0;
wire R10C28_X01;
wire R20C31_GB30;
wire R10C7_B2;
wire R21C35_GB00;
wire R28C28_N25;
wire R10C29_F5;
wire R4C21_GB30;
wire R1C47_D2;
wire R5C8_GB30;
wire R8C15_GB10;
wire R10C28_D1;
wire R21C25_GB20;
wire R3C9_GB50;
wire R14C23_GB50;
wire R7C46_GB40;
wire R21C29_GT10;
wire R2C42_GT00;
wire R11C46_GB50;
wire R4C33_GB70;
wire R1C1_CLK1;
wire R28C46_S81;
wire R11C25_GT10;
wire R20C23_SPINE17;
wire R23C36_GT00;
wire R15C42_GT00;
wire R28C43_N23;
wire R1C28_E12;
wire R21C5_GB00;
wire R17C9_GB40;
wire R2C25_GB60;
wire R25C5_GBO0;
wire R12C42_GB20;
wire R16C12_GBO0;
wire R20C6_GB70;
wire R13C13_GB60;
wire R17C22_GB50;
wire R9C32_GT10;
wire R21C15_GB70;
wire R5C37_GB50;
wire R13C28_GB60;
wire R10C37_E80;
wire R10C40_SEL3;
wire R4C8_GT10;
wire R28C37_Q2;
wire R18C5_GB40;
wire R10C30_N24;
wire R28C28_Q3;
wire R5C25_GB10;
wire R23C22_GBO0;
wire R16C31_GB60;
wire R25C26_GB50;
wire R27C43_GT10;
wire R15C30_GBO0;
wire R25C46_GB40;
wire R16C23_GB00;
wire R5C20_GB10;
wire R24C18_GBO1;
wire R11C35_GB70;
wire R10C30_LSR1;
wire R17C46_GB30;
wire R11C18_GBO0;
wire R23C25_GB30;
wire R8C30_GB20;
wire R14C37_GB30;
wire R5C20_GB30;
wire R8C32_GT00;
wire R28C4_E12;
wire R22C3_GB70;
wire R6C42_GT00;
wire R21C24_GB60;
wire R26C33_GB10;
wire R6C33_GB30;
wire R10C7_C6;
wire R2C42_GB70;
wire R15C17_GB10;
wire R6C34_GT00;
wire R13C33_GB60;
wire R3C9_GBO0;
wire R10C26_N81;
wire R28C46_CE2;
wire R26C14_GT10;
wire R28C4_X03;
wire R3C39_GB70;
wire R15C10_GB10;
wire R15C40_GB30;
wire R8C22_GB40;
wire R18C10_GT10;
wire R15C10_GB70;
wire R17C10_GB10;
wire R17C44_GB70;
wire R25C16_GB30;
wire R10C30_E22;
wire R28C40_A4;
wire R3C31_GB60;
wire R21C29_GB60;
wire R13C7_GB30;
wire R28C31_SEL4;
wire R21C25_GB40;
wire R20C45_GB30;
wire R28C7_Q4;
wire R18C27_GB40;
wire R3C30_GB10;
wire R28C7_SEL1;
wire R9C3_GBO0;
wire R27C26_GB00;
wire R17C8_GB00;
wire R17C46_GBO0;
wire R24C38_GT00;
wire R10C31_SN10;
wire R28C19_N81;
wire R29C28_A2;
wire R25C45_GBO1;
wire R10C13_S24;
wire R14C25_GB60;
wire R2C33_GB20;
wire R10C43_W20;
wire R7C10_GT10;
wire R9C44_GB40;
wire R23C34_GB00;
wire R28C37_S83;
wire R8C28_GB10;
wire R20C2_GB20;
wire R14C43_GB70;
wire R17C42_GT10;
wire R16C33_GB10;
wire R10C19_F2;
wire R28C40_C7;
wire R28C13_S13;
wire R10C10_B3;
wire R10C13_E21;
wire R28C37_N82;
wire R28C7_A6;
wire R16C11_GB30;
wire R10C10_W22;
wire R26C6_GB00;
wire R16C43_GT00;
wire R28C19_W20;
wire R24C6_GB30;
wire R18C18_GT00;
wire R13C17_GB30;
wire R20C26_GT00;
wire R20C36_GT00;
wire R10C30_E13;
wire R12C38_GB50;
wire R5C15_GT10;
wire R13C29_GBO1;
wire R27C4_GT00;
wire R15C2_GB50;
wire R2C10_GB30;
wire R10C29_LSR2;
wire R6C40_GB70;
wire R28C19_D5;
wire R14C40_GBO1;
wire R22C46_GBO0;
wire R5C39_GB30;
wire R28C28_S23;
wire R10C31_E21;
wire R3C44_GT00;
wire R22C7_GB40;
wire R17C3_GB30;
wire R20C41_GB10;
wire R25C30_GB70;
wire R16C42_GB40;
wire R23C27_GB30;
wire R6C38_GBO0;
wire R14C37_GT10;
wire R12C26_GB30;
wire R10C16_E24;
wire R13C22_GB30;
wire R26C11_GB40;
wire R4C21_GB40;
wire R14C10_GT00;
wire R24C41_GBO0;
wire R10C30_S81;
wire R5C21_GB10;
wire R17C31_GB10;
wire R10C22_B7;
wire R6C21_GB00;
wire R27C30_GB30;
wire R17C22_GT10;
wire R24C34_GB10;
wire R23C38_GT10;
wire R13C11_GB00;
wire R10C31_N82;
wire R18C45_GB40;
wire R21C16_GBO0;
wire R28C31_S22;
wire R5C46_GB40;
wire R10C26_X06;
wire R25C43_GT00;
wire R10C43_W10;
wire R9C45_GBO0;
wire R5C12_GB00;
wire R10C31_W26;
wire R12C4_GB50;
wire R22C24_GB70;
wire R12C46_GB00;
wire R4C6_GBO0;
wire R10C30_S11;
wire R11C21_GB00;
wire R10C25_N81;
wire R28C13_SEL1;
wire R26C3_GB10;
wire R18C24_GB20;
wire R6C5_GBO0;
wire R16C8_GBO1;
wire R11C18_GB70;
wire R11C31_GBO0;
wire R28C31_D6;
wire R9C3_GBO1;
wire R15C9_GT10;
wire R10C10_N25;
wire R25C40_GB20;
wire R26C16_GB10;
wire R17C18_GB50;
wire R23C3_GB70;
wire R3C45_GB20;
wire R6C31_GB50;
wire R17C26_GB60;
wire R10C22_S20;
wire R28C4_Q5;
wire R23C20_GB00;
wire R10C28_C1;
wire R22C34_GT00;
wire R26C7_GB20;
wire R26C7_GB00;
wire R2C21_GB20;
wire R2C25_GT00;
wire R20C18_GBO0;
wire R28C13_C1;
wire R28C13_N13;
wire R28C31_B7;
wire R11C34_GT10;
wire R23C38_GT00;
wire R27C9_GBO0;
wire R6C13_GT00;
wire R5C31_GB40;
wire R11C2_GB60;
wire R28C37_E10;
wire R24C24_GB50;
wire R8C12_GB30;
wire R6C23_GB30;
wire R13C11_GB20;
wire R13C16_GB50;
wire R26C26_GB70;
wire R9C34_GBO1;
wire R10C16_A0;
wire R7C44_GB00;
wire R9C36_GB30;
wire R10C26_C6;
wire R13C38_GBO1;
wire R28C28_B5;
wire R6C42_GBO1;
wire R22C36_GB20;
wire R25C13_GB30;
wire R10C16_S25;
wire R6C1_GT00;
wire R14C15_GB60;
wire R28C28_B7;
wire R16C19_GB40;
wire R6C13_GBO0;
wire R17C6_GB50;
wire R2C41_GB60;
wire R12C41_GBO1;
wire R22C19_GBO1;
wire R5C39_GBO1;
wire R10C22_E21;
wire R28C19_D7;
wire R2C36_SPINE0;
wire R2C4_GT10;
wire R17C44_GB10;
wire R12C3_GBO0;
wire R12C31_GBO1;
wire R2C6_GB50;
wire R1C32_D1;
wire R26C30_GB60;
wire R11C37_GB10;
wire R20C17_GB20;
wire R2C37_GT00;
wire R18C45_GB10;
wire R21C7_GT00;
wire R6C36_GT00;
wire R10C27_X01;
wire R10C30_W20;
wire R28C25_N20;
wire R24C35_GB40;
wire R9C15_GT00;
wire R8C5_GBO0;
wire R2C15_GBO1;
wire R25C36_GB40;
wire R11C5_GB30;
wire R28C28_C3;
wire R8C29_GB40;
wire R4C46_GT00;
wire R20C8_SPINE20;
wire R21C46_GB10;
wire R1C1_E22;
wire R15C5_GB60;
wire R10C10_S22;
wire R29C28_S22;
wire R3C24_GB00;
wire R14C25_GB30;
wire R10C26_A0;
wire R3C26_GT10;
wire R28C7_F1;
wire R22C16_GB50;
wire R28C34_C1;
wire R12C36_GB50;
wire R29C28_F0;
wire R28C13_X06;
wire R2C12_GB00;
wire R22C21_GB30;
wire R25C34_GBO1;
wire R17C7_GB70;
wire R27C12_GT10;
wire R1C1_D4;
wire R12C18_GT10;
wire R21C18_GB00;
wire R22C27_GB10;
wire R16C18_GB30;
wire R7C35_GB10;
wire R8C16_GB10;
wire R1C47_SEL2;
wire R4C42_GB30;
wire R6C45_GBO0;
wire R1C28_SEL2;
wire R4C22_GB70;
wire R28C10_D1;
wire R12C45_GB60;
wire R27C1_GBO1;
wire R28C22_S81;
wire R11C20_GB60;
wire R14C23_GB70;
wire R2C14_GB40;
wire R9C13_GB40;
wire R17C3_GBO1;
wire R28C31_C0;
wire R21C19_GBO1;
wire R9C32_GB70;
wire R17C16_GT10;
wire R6C45_GT10;
wire R1C32_E23;
wire R15C22_GB20;
wire R1C32_CLK1;
wire R14C31_GB70;
wire R24C29_GB60;
wire R5C5_GB30;
wire R6C11_GB70;
wire R5C5_GB00;
wire R10C30_E83;
wire R28C19_CE0;
wire R14C40_GB10;
wire R3C5_GB70;
wire R11C9_GB30;
wire R1C47_LSR2;
wire R4C10_GBO1;
wire R10C40_S80;
wire R21C29_GBO0;
wire R8C26_GB40;
wire R11C19_GBO0;
wire R5C46_GBO1;
wire R1C1_S23;
wire R10C29_S10;
wire R9C33_GB70;
wire R17C22_GB10;
wire R28C37_X04;
wire R9C19_GB30;
wire R10C16_SEL1;
wire R6C13_GT10;
wire R27C20_GBO1;
wire R16C36_GB70;
wire R28C43_D4;
wire R10C28_W82;
wire R9C4_GBO1;
wire R16C26_GBO0;
wire R27C36_GB00;
wire R8C2_GB50;
wire R13C34_GB50;
wire R16C8_GB40;
wire R12C39_GB70;
wire R20C46_GT10;
wire R28C37_SEL5;
wire R10C43_N82;
wire R22C29_GB30;
wire R10C26_F0;
wire R10C29_Q4;
wire R10C10_CE0;
wire R10C37_B2;
wire R4C39_GB60;
wire R25C11_GT00;
wire R4C27_GBO0;
wire R10C28_S12;
wire R24C43_GB60;
wire R2C21_GT00;
wire R20C5_GB20;
wire R4C36_GBO0;
wire R27C32_GT00;
wire R10C7_F2;
wire R8C26_GB10;
wire R12C29_GB60;
wire R25C4_GT10;
wire R1C1_Q3;
wire R13C34_GB60;
wire R27C6_GBO0;
wire R12C16_GB50;
wire R18C45_GB60;
wire R3C11_GB40;
wire R22C14_GBO1;
wire R6C42_GB50;
wire R5C30_GBO0;
wire R2C15_GB50;
wire R1C1_W23;
wire R10C37_Q4;
wire R2C16_GB10;
wire R28C22_S12;
wire R23C26_GB30;
wire R6C10_GBO1;
wire R15C8_GB20;
wire R10C25_A6;
wire R28C40_LSR1;
wire R6C23_GBO0;
wire R5C1_GBO0;
wire R18C4_GBO0;
wire R10C13_A3;
wire R8C11_GB40;
wire R14C22_GB50;
wire R26C20_GB70;
wire R10C7_S82;
wire R28C22_F5;
wire R28C34_E82;
wire R21C41_GBO1;
wire R13C22_GBO0;
wire R1C32_B7;
wire R23C16_GB10;
wire R11C21_GB10;
wire R10C7_E80;
wire R10C34_B5;
wire R28C10_S81;
wire R20C22_GB20;
wire R2C41_SPINE3;
wire R5C6_GB40;
wire R13C10_GBO1;
wire R20C3_GBO1;
wire R7C39_GB40;
wire R11C37_GB70;
wire R8C32_GB50;
wire R8C46_GB70;
wire R26C35_GB30;
wire R18C40_GB70;
wire R15C12_GB10;
wire R14C9_GB30;
wire R15C3_GB20;
wire R24C8_GB20;
wire R4C9_GB60;
wire R22C27_GB40;
wire R4C12_GB40;
wire R9C3_GB20;
wire R27C26_GB10;
wire R23C40_GB60;
wire R1C28_X03;
wire R15C45_GB40;
wire R10C34_E13;
wire R26C36_GB30;
wire R28C43_N27;
wire R18C13_GBO1;
wire R2C1_GT10;
wire R4C13_GB70;
wire R24C23_GBO0;
wire R20C14_SPINE18;
wire R18C4_GB70;
wire R28C40_F2;
wire R22C28_GB30;
wire R14C44_GB30;
wire R25C42_GBO0;
wire R10C10_W21;
wire R22C43_GT10;
wire R16C6_GT00;
wire R4C21_GBO1;
wire R24C17_GBO0;
wire R12C42_GB40;
wire R7C22_GT00;
wire R28C40_F5;
wire R23C9_GB50;
wire R15C37_GB40;
wire R14C6_GBO1;
wire R7C25_GBO0;
wire R8C37_GB70;
wire R6C29_GT10;
wire R13C46_GBO1;
wire R28C31_S11;
wire R4C10_GB70;
wire R15C7_GB10;
wire R10C27_D4;
wire R28C22_E11;
wire R25C5_GT00;
wire R13C39_GB00;
wire R5C43_GB10;
wire R1C28_S24;
wire R16C14_GB70;
wire R10C31_N83;
wire R25C11_GB30;
wire R25C34_GB60;
wire R10C30_E80;
wire R28C28_LSR0;
wire R26C29_GBO0;
wire R18C45_GB50;
wire R28C28_E82;
wire R6C46_GB40;
wire R14C12_GB10;
wire R3C29_GB10;
wire R16C42_GB70;
wire R24C11_GB10;
wire R2C26_GB50;
wire R1C32_S80;
wire R28C10_SEL2;
wire R2C7_SPINE9;
wire R5C8_GBO0;
wire R10C31_E82;
wire R18C31_GB10;
wire R18C4_GT10;
wire R7C42_GBO0;
wire R10C43_Q0;
wire R15C19_GBO1;
wire R10C40_Q5;
wire R25C13_GB20;
wire R25C10_GT10;
wire R2C13_GBO1;
wire R18C17_GBO1;
wire R27C23_GBO1;
wire R6C4_GB00;
wire R4C4_GB20;
wire R5C17_GB20;
wire R16C3_GT10;
wire R14C28_GB40;
wire R9C37_GB10;
wire R23C44_GB60;
wire R21C43_GT00;
wire R28C28_E21;
wire R15C41_GB50;
wire R20C24_GB10;
wire R7C19_GB70;
wire R7C2_GB60;
wire R22C8_GBO0;
wire R2C5_GB30;
wire R20C5_GB50;
wire R27C33_GB70;
wire R15C42_GB70;
wire R10C30_SPINE3;
wire R28C13_F6;
wire R28C4_W25;
wire R1C1_S13;
wire R28C31_LSR1;
wire R20C7_GBO1;
wire R18C3_GT00;
wire R11C3_GBO0;
wire R26C32_GB50;
wire R15C41_GB10;
wire R16C45_GB50;
wire R22C10_GB30;
wire R23C13_GB20;
wire R7C13_GBO0;
wire R20C36_SPINE28;
wire R28C46_D3;
wire R6C27_GB50;
wire R5C29_GB30;
wire R10C27_N10;
wire R28C10_SN10;
wire R23C27_GB40;
wire R13C44_GB00;
wire R11C22_GB00;
wire R22C25_GB50;
wire R23C17_GB60;
wire R10C13_SEL2;
wire R8C12_GT10;
wire R1C1_S12;
wire R16C37_GT00;
wire R1C28_SEL4;
wire R2C3_GB00;
wire R28C22_X08;
wire R28C34_F6;
wire R12C23_GB10;
wire R28C7_X02;
wire R20C29_GB00;
wire R21C42_GBO1;
wire R10C16_Q0;
wire R5C21_GB30;
wire R3C15_GB50;
wire R28C16_N21;
wire R10C13_SEL1;
wire R28C37_B7;
wire R20C5_GB10;
wire R8C11_GB10;
wire R14C7_GB20;
wire R26C3_GB00;
wire R9C4_GB70;
wire R18C31_GB20;
wire R20C3_GB00;
wire R16C19_GB50;
wire R28C4_W13;
wire R6C18_GBO1;
wire R23C36_GBO1;
wire R11C45_GB10;
wire R15C16_GB20;
wire R12C18_GB00;
wire R10C29_W11;
wire R24C32_GB40;
wire R11C36_GB50;
wire R10C43_N11;
wire R17C27_GT10;
wire R15C6_GT10;
wire R18C44_GB10;
wire R28C28_B6;
wire R25C16_GB50;
wire R10C40_E13;
wire R28C43_E22;
wire R18C14_GB30;
wire R13C40_GB40;
wire R18C18_GBO0;
wire R28C31_X03;
wire R23C7_GT00;
wire R10C27_W10;
wire R14C2_GB30;
wire R21C11_GB70;
wire R26C23_GB10;
wire R12C25_GBO0;
wire R26C6_GB70;
wire R10C40_W12;
wire R10C10_S25;
wire R22C30_GB60;
wire R10C31_C2;
wire R6C20_GT10;
wire R28C16_C7;
wire R28C43_CLK2;
wire R28C37_D7;
wire R20C17_GBO1;
wire R23C5_GB70;
wire R28C16_W20;
wire R3C4_GB10;
wire R6C40_GT10;
wire R24C39_GT00;
wire R25C15_GB10;
wire R8C3_GB40;
wire R28C16_F4;
wire R7C39_GBO0;
wire R10C25_C6;
wire R7C23_GT10;
wire R17C26_GB40;
wire R2C27_SPINE9;
wire R9C45_GT00;
wire R7C27_GBO0;
wire R10C13_W25;
wire R18C9_GB20;
wire R26C42_GBO0;
wire R28C4_E20;
wire R28C43_D2;
wire R28C10_X08;
wire R5C31_GT10;
wire R28C40_C5;
wire R2C32_GBO0;
wire R10C27_S81;
wire R12C26_GT10;
wire R23C6_GB30;
wire R27C7_GB50;
wire R28C16_A0;
wire R4C24_GB70;
wire R13C17_GB10;
wire R21C36_GT00;
wire R10C37_W81;
wire R6C9_GB00;
wire R28C43_Q1;
wire R28C22_F0;
wire R5C41_GT00;
wire R21C45_GB00;
wire R3C23_GB50;
wire R22C6_GBO0;
wire R26C25_GB70;
wire R10C22_F1;
wire R11C22_GBO0;
wire R10C30_Q5;
wire R12C4_GB60;
wire R10C40_A5;
wire R6C32_GT10;
wire R6C43_GBO0;
wire R20C28_GT10;
wire R2C20_GB00;
wire R26C28_GB00;
wire R14C44_GB20;
wire R9C37_GT10;
wire R4C18_GB30;
wire R27C43_GB40;
wire R20C44_GB00;
wire R21C6_GT10;
wire R13C25_GT00;
wire R2C25_GB00;
wire R7C11_GB10;
wire R7C14_GB70;
wire R16C40_GB10;
wire R6C44_GB40;
wire R15C44_GB30;
wire R23C26_GB00;
wire R28C37_SEL7;
wire R3C10_GB60;
wire R5C35_GT10;
wire R16C14_GB20;
wire R7C34_GB30;
wire R12C30_GBO0;
wire R20C36_GB20;
wire R15C36_GB60;
wire R10C28_Q3;
wire R13C12_GB00;
wire R3C33_GBO1;
wire R2C32_GB30;
wire R10C22_N11;
wire R10C34_W13;
wire R14C4_GB30;
wire R18C16_GB60;
wire R11C9_GBO0;
wire R23C24_GB60;
wire R2C44_GB70;
wire R1C28_F1;
wire R17C12_GB30;
wire R2C6_GB40;
wire R9C40_GB20;
wire R3C7_GB10;
wire R28C13_W83;
wire R10C29_F4;
wire R28C31_W12;
wire R14C35_GT10;
wire R15C39_GB20;
wire R20C18_GB20;
wire R21C14_GB20;
wire R18C9_GB00;
wire R18C37_GB30;
wire R16C14_GB10;
wire R12C37_GBO0;
wire R9C3_GB30;
wire R23C24_GB70;
wire R13C17_GB60;
wire R2C34_GB70;
wire R3C3_GBO1;
wire R11C35_GB40;
wire R17C10_GT10;
wire R26C9_GT00;
wire R1C28_Q5;
wire R10C16_W81;
wire R28C25_N11;
wire R3C26_GBO0;
wire R28C37_N10;
wire R5C11_GT00;
wire R25C34_GT00;
wire R27C45_GBO0;
wire R10C13_E13;
wire R4C25_GB10;
wire R7C4_GB50;
wire R2C4_GB30;
wire R10C31_F4;
wire R22C37_GB50;
wire R6C23_GT00;
wire R10C43_E11;
wire R28C40_E26;
wire R14C21_GB20;
wire R25C6_GT00;
wire R1C32_S23;
wire R2C35_GB00;
wire R26C27_GT10;
wire R22C1_GT00;
wire R7C3_GBO0;
wire R10C13_C0;
wire R10C29_CE2;
wire R21C2_GT10;
wire R9C19_GB60;
wire R10C40_F2;
wire R9C20_GB20;
wire R9C9_GT00;
wire R8C35_GB10;
wire R6C28_GB70;
wire R28C22_N21;
wire R3C23_GT10;
wire R23C40_GT00;
wire R9C12_GB50;
wire R14C19_GBO0;
wire R23C37_GB40;
wire R15C13_GB40;
wire R15C20_GB60;
wire R10C16_E11;
wire R28C4_EW20;
wire R8C18_GB70;
wire R15C34_GB40;
wire R23C18_GT00;
wire R18C26_GB00;
wire R14C9_GB40;
wire R5C40_GB30;
wire R7C6_GBO1;
wire R2C33_GT00;
wire R3C22_GB30;
wire R11C29_GB40;
wire R8C9_GBO1;
wire R9C4_GB30;
wire R10C25_W20;
wire R24C27_GBO0;
wire R6C11_GB50;
wire R28C10_CLK1;
wire R16C39_GB20;
wire R7C40_GB10;
wire R6C35_GB30;
wire R3C43_GB50;
wire R12C32_GB60;
wire R20C19_GB40;
wire R15C33_GB30;
wire R10C26_A4;
wire R10C25_E13;
wire R17C2_GB10;
wire R10C43_E20;
wire R21C42_GB00;
wire R24C25_GB40;
wire R12C37_GB30;
wire R8C13_GB70;
wire R23C7_GB70;
wire R12C38_GT00;
wire R25C25_GB30;
wire R8C45_GB10;
wire R28C46_E25;
wire R17C2_GT10;
wire R7C9_GB20;
wire R13C31_GB70;
wire R15C39_GB70;
wire R23C36_GB70;
wire R15C40_GT00;
wire R11C32_GT00;
wire R24C6_GB60;
wire R10C22_W20;
wire R10C34_Q1;
wire R28C19_E80;
wire R12C7_GT10;
wire R15C2_GB30;
wire R17C30_GT00;
wire R20C40_GBO0;
wire R24C31_GT10;
wire R27C16_GB00;
wire R4C24_GBO0;
wire R9C27_GB20;
wire R12C8_GB30;
wire R16C14_GB30;
wire R23C10_GB50;
wire R26C13_GB60;
wire R18C28_GT10;
wire R27C26_GB20;
wire R3C38_GB60;
wire R15C24_GT00;
wire R10C25_N25;
wire R12C42_GB70;
wire R11C21_GB60;
wire R21C36_GB10;
wire R24C46_GB00;
wire R6C24_GB60;
wire R14C42_GB60;
wire R10C29_SN10;
wire R10C31_S21;
wire R8C12_GB70;
wire R28C10_A3;
wire R16C10_GT10;
wire R18C12_GB30;
wire R28C37_N26;
wire R15C31_GB00;
wire R14C24_GB30;
wire R10C26_N10;
wire R28C28_N21;
wire R15C24_GB40;
wire R6C42_GB20;
wire R7C23_GB30;
wire R12C28_GB10;
wire R27C32_GB30;
wire R1C28_N23;
wire R10C22_N24;
wire R10C26_S81;
wire R20C7_GB40;
wire R28C43_C5;
wire R16C27_GB50;
wire R10C28_Q1;
wire R8C18_GB30;
wire R12C7_GB00;
wire R13C34_GBO0;
wire R1C1_S81;
wire R4C19_GB60;
wire R11C32_GB40;
wire R1C1_N20;
wire R20C21_GB70;
wire R13C22_GBO1;
wire R10C25_D0;
wire R22C12_GB10;
wire R25C24_GB40;
wire R6C21_GB20;
wire R12C40_GB40;
wire R7C16_GBO0;
wire R1C1_D2;
wire R28C4_W22;
wire R10C43_N12;
wire R28C28_S25;
wire R5C10_GT00;
wire R22C6_GB60;
wire R21C34_GBO0;
wire R10C16_SEL6;
wire R7C32_GB30;
wire R12C37_GB10;
wire R10C28_N21;
wire R16C39_GB60;
wire R27C14_GB60;
wire R4C30_GB00;
wire R11C15_GT00;
wire R6C10_GB10;
wire R13C39_GBO1;
wire R23C30_GB00;
wire R10C27_W24;
wire R13C25_GB60;
wire R7C36_GB20;
wire R25C4_GT00;
wire R3C16_GB00;
wire R15C46_GB50;
wire R10C34_A3;
wire R9C12_GB10;
wire R7C20_GB50;
wire R4C43_GB50;
wire R6C43_GT00;
wire R18C26_GB40;
wire R28C13_N21;
wire R10C19_W25;
wire R20C43_GB30;
wire R10C27_SPINE13;
wire R14C42_GB20;
wire R7C41_GT10;
wire R10C26_C2;
wire R28C16_W13;
wire R25C40_GB10;
wire R26C18_GBO0;
wire R28C7_E26;
wire R17C14_GT10;
wire R4C21_GB50;
wire R20C10_GB70;
wire R10C22_N10;
wire R13C37_GB10;
wire R10C29_Q3;
wire R21C34_GB70;
wire R29C28_A0;
wire R10C37_W83;
wire R16C9_GB10;
wire R13C44_GT10;
wire R10C37_W22;
wire R28C19_F2;
wire R6C23_GB20;
wire R18C34_GBO0;
wire R28C25_S22;
wire R12C32_GBO1;
wire R17C24_GB10;
wire R21C46_GB70;
wire R10C10_SN10;
wire R4C37_GT00;
wire R6C2_GT00;
wire R28C46_W13;
wire R10C25_E20;
wire R20C40_GB50;
wire R10C30_N23;
wire R16C7_GBO1;
wire R12C1_GT10;
wire R24C45_GB60;
wire R2C16_GT10;
wire R14C29_GT10;
wire R5C33_GB20;
wire R9C2_GT10;
wire R16C34_GB40;
wire R1C28_W82;
wire R10C30_N13;
wire R6C18_GB60;
wire R10C7_A2;
wire R23C2_GBO0;
wire R12C41_GB40;
wire R28C43_N11;
wire R29C28_W10;
wire R17C45_GT00;
wire R13C46_GB00;
wire R9C31_GB10;
wire R1C28_S10;
wire R10C27_SPINE10;
wire R18C25_GT00;
wire R3C39_GB40;
wire R15C5_GB50;
wire R23C32_GB10;
wire R28C19_E22;
wire R25C38_GT00;
wire R2C17_GB60;
wire R21C14_GT00;
wire R27C38_GB70;
wire R13C2_GBO1;
wire R28C43_A4;
wire R11C42_GBO1;
wire R4C26_GT00;
wire R23C42_GBO0;
wire R22C28_GB20;
wire R10C27_SEL2;
wire R28C25_D2;
wire R4C3_GB20;
wire R25C32_GT10;
wire R17C8_GB70;
wire R10C7_S11;
wire R10C43_A6;
wire R6C21_GB30;
wire R11C10_GB50;
wire R7C25_GB50;
wire R25C43_GT10;
wire R10C25_W12;
wire R10C30_B0;
wire R17C8_GB60;
wire R11C16_GB70;
wire R23C17_GB70;
wire R8C8_GBO0;
wire R28C10_D7;
wire R1C28_S22;
wire R1C1_SEL7;
wire R14C8_GB40;
wire R16C19_GT10;
wire R16C7_GB50;
wire R20C13_GBO1;
wire R24C44_GB40;
wire R12C10_GT00;
wire R5C43_GB30;
wire R25C29_GB50;
wire R7C11_GT00;
wire R22C46_GB00;
wire R6C17_GT10;
wire R13C39_GT00;
wire R2C18_GB10;
wire R10C25_SN10;
wire R10C29_D1;
wire R29C28_SEL5;
wire R15C25_GB60;
wire R11C32_GB70;
wire R28C7_D7;
wire R10C13_B4;
wire R12C5_GT10;
wire R17C30_GB10;
wire R28C10_W26;
wire R14C11_GB40;
wire R10C16_CE2;
wire R17C23_GB60;
wire R21C18_GBO1;
wire R6C40_GB00;
wire R21C33_GB10;
wire R18C25_GB60;
wire R24C18_GB70;
wire R7C30_GB20;
wire R17C42_GB60;
wire R26C5_GB60;
wire R27C32_GB00;
wire R5C6_GB60;
wire R25C14_GB40;
wire R1C32_S83;
wire R28C13_W26;
wire R13C21_GBO1;
wire R4C20_GB30;
wire R8C33_GB70;
wire R7C27_GT00;
wire R2C26_GBO1;
wire R20C35_SPINE29;
wire R27C39_GT00;
wire R18C38_GB40;
wire R23C44_GBO0;
wire R10C31_F7;
wire R11C15_GBO0;
wire R5C37_GT10;
wire R24C38_GT10;
wire R21C16_GB70;
wire R10C40_F6;
wire R11C28_GB60;
wire R28C28_SEL2;
wire R9C31_GBO0;
wire R17C34_GBO0;
wire R7C5_GB00;
wire R23C18_GB70;
wire R20C14_GB70;
wire R27C15_GB30;
wire R27C39_GB70;
wire R4C34_GB60;
wire R10C43_EW20;
wire R12C21_GBO1;
wire R9C17_GB50;
wire R17C10_GB60;
wire R14C28_GT10;
wire R8C1_GBO1;
wire R20C11_GT10;
wire R14C8_GB50;
wire R10C29_LSR0;
wire R2C30_GB50;
wire R28C34_D7;
wire R2C37_GB20;
wire R10C37_B7;
wire R6C34_GB30;
wire R17C15_GB40;
wire R25C29_GB20;
wire R8C40_GB10;
wire R23C6_GB20;
wire R10C22_S23;
wire R9C3_GB70;
wire R15C27_GBO0;
wire R10C27_F7;
wire R28C19_Q7;
wire R9C2_GT00;
wire R26C6_GBO1;
wire R25C30_GBO0;
wire R10C26_B2;
wire R26C43_GB60;
wire R11C22_GB70;
wire R28C10_S13;
wire R28C7_D3;
wire R16C7_GB20;
wire R28C16_SN10;
wire R28C43_Q3;
wire R28C28_F2;
wire R22C16_GB30;
wire R3C36_GB50;
wire R18C32_GT00;
wire R6C12_GB70;
wire R18C2_GB20;
wire R5C7_GB00;
wire R10C22_N82;
wire R10C28_B0;
wire R9C35_GBO1;
wire R27C2_GB40;
wire R12C23_GB00;
wire R26C13_GB70;
wire R10C10_E23;
wire R6C14_GB70;
wire R4C31_GB40;
wire R16C1_GBO1;
wire R20C6_GBO0;
wire R10C31_E26;
wire R28C34_X03;
wire R3C7_GT10;
wire R18C17_GB40;
wire R16C27_GB60;
wire R17C39_GB60;
wire R20C44_SPINE28;
wire R25C5_GB10;
wire R24C17_GT00;
wire R24C2_GT00;
wire R9C41_GB50;
wire R8C31_GBO1;
wire R18C35_GB10;
wire R16C46_GT00;
wire R26C31_GB40;
wire R15C4_GB10;
wire R16C44_GB60;
wire R24C14_GB60;
wire R1C28_S80;
wire R8C46_GB20;
wire R5C40_GB00;
wire R3C13_GB70;
wire R20C19_GB10;
wire R5C30_GBO1;
wire R13C39_GB40;
wire R18C31_GB70;
wire R10C10_C1;
wire R14C23_GT10;
wire R13C27_GB00;
wire R20C5_GB60;
wire R12C34_GBO0;
wire R25C30_GT10;
wire R2C7_GBO1;
wire R28C7_SEL0;
wire R21C26_GT10;
wire R25C16_GBO1;
wire R22C36_GB60;
wire R28C43_E26;
wire R20C46_GB50;
wire R17C25_GB50;
wire R10C27_N21;
wire R28C46_Q2;
wire R11C16_GB20;
wire R12C5_GT00;
wire R14C45_GBO0;
wire R1C47_SEL3;
wire R13C14_GT10;
wire R28C25_B5;
wire R5C16_GB30;
wire R13C7_GBO0;
wire R25C28_GB70;
wire R23C1_GT10;
wire R10C30_S25;
wire R16C25_GT10;
wire R10C30_X06;
wire R28C46_S24;
wire R23C26_GBO0;
wire R10C30_D2;
wire R18C36_GB70;
wire R1C1_N11;
wire R10C43_E82;
wire R28C31_C5;
wire R29C28_C1;
wire R13C32_GBO0;
wire R10C19_CE0;
wire R5C19_GB70;
wire R22C23_GB10;
wire R15C11_GB70;
wire R10C16_SEL5;
wire R28C19_S26;
wire R10C28_A2;
wire R22C5_GT00;
wire R22C1_GBO1;
wire R7C30_GBO0;
wire R13C5_GT00;
wire R10C27_N80;
wire R8C36_GT10;
wire R10C37_N82;
wire R9C18_GB20;
wire R10C22_E80;
wire R10C40_N25;
wire R28C16_W80;
wire R28C43_CE1;
wire R17C17_GB60;
wire R5C4_GBO0;
wire R25C42_GB10;
wire R27C44_GB40;
wire R14C29_GB30;
wire R10C31_E11;
wire R22C40_GB30;
wire R10C25_E80;
wire R14C19_GT00;
wire R6C17_GB30;
wire R28C25_N82;
wire R8C8_GT10;
wire R8C3_GBO1;
wire R2C46_GBO1;
wire R20C34_SPINE26;
wire R28C25_B2;
wire R14C32_GB20;
wire R27C29_GB10;
wire R26C2_GB20;
wire R18C34_GT00;
wire R28C37_N83;
wire R27C5_GB40;
wire R3C4_GBO1;
wire R20C27_SPINE17;
wire R2C34_GB60;
wire R1C32_D6;
wire R21C46_GT10;
wire R10C7_N25;
wire R23C29_GB20;
wire R15C46_GB40;
wire R10C37_D0;
wire R10C29_F0;
wire R16C27_GB70;
wire R16C43_GB30;
wire R10C43_SN10;
wire R2C3_GB50;
wire R13C29_GBO0;
wire R18C31_GB60;
wire R7C24_GBO0;
wire R28C28_E22;
wire R29C28_N26;
wire R6C3_GT10;
wire R8C30_GB00;
wire R9C38_GB40;
wire R1C28_A7;
wire R10C28_UNK125;
wire R14C17_GB10;
wire R28C13_E12;
wire R26C9_GT10;
wire R18C2_GB00;
wire R14C44_GB40;
wire R15C12_GBO1;
wire R10C40_E22;
wire R21C39_GB10;
wire R10C26_N23;
wire R18C44_GB60;
wire R10C26_W82;
wire R10C19_D3;
wire R21C30_GB50;
wire R14C18_GB60;
wire R24C24_GB40;
wire R5C24_GB50;
wire R16C20_GT10;
wire R5C2_GB50;
wire R13C12_GBO0;
wire R5C23_GB60;
wire R18C27_GB70;
wire R17C22_GBO0;
wire R28C4_N80;
wire R2C37_GB00;
wire R20C41_SPINE27;
wire R9C12_GBO1;
wire R2C8_SPINE8;
wire R12C33_GB30;
wire R5C24_GB20;
wire R7C36_GT00;
wire R11C39_GT00;
wire R25C16_GB40;
wire R13C36_GB00;
wire R3C34_GB30;
wire R26C31_GB60;
wire R28C16_X08;
wire R10C22_E83;
wire R24C32_GT10;
wire R25C1_GT10;
wire R6C44_GB00;
wire R10C13_N23;
wire R27C4_GT10;
wire R4C31_GB00;
wire R24C24_GB20;
wire R21C3_GT00;
wire R27C41_GB50;
wire R10C13_W24;
wire R9C38_GB50;
wire R2C4_GT00;
wire R14C39_GB50;
wire R8C29_GT00;
wire R11C26_GT10;
wire R18C12_GB00;
wire R8C2_GB70;
wire R2C9_GB60;
wire R25C27_GB50;
wire R13C4_GB60;
wire R15C6_GBO0;
wire R6C26_GT10;
wire R10C13_F5;
wire R2C34_GB10;
wire R3C16_GT10;
wire R28C46_Q3;
wire R18C19_GB00;
wire R10C31_N12;
wire R28C16_C6;
wire R27C40_GT00;
wire R2C14_GB70;
wire R20C4_GB20;
wire R9C34_GB30;
wire R7C40_GB70;
wire R28C19_Q5;
wire R10C43_D5;
wire R24C36_GB50;
wire R10C10_D4;
wire R14C24_GB50;
wire R20C37_GB40;
wire R1C47_W20;
wire R13C42_GB30;
wire R6C4_GB30;
wire R28C4_X06;
wire R23C27_GT00;
wire R26C40_GB60;
wire R10C22_N81;
wire R3C2_GT10;
wire R2C35_GB10;
wire R28C34_W82;
wire R28C13_S10;
wire R13C32_GB60;
wire R1C1_A3;
wire R5C44_GB50;
wire R10C22_Q0;
wire R7C16_GB60;
wire R2C8_GB20;
wire R6C31_GB30;
wire R10C31_SEL5;
wire R28C28_S82;
wire R28C28_X05;
wire R28C37_E27;
wire R28C46_F6;
wire R16C17_GBO1;
wire R23C38_GB50;
wire R20C35_GBO0;
wire R28C25_W27;
wire R28C28_CLK1;
wire R11C3_GT10;
wire R13C37_GB40;
wire R20C9_GB50;
wire R28C28_SEL1;
wire R4C24_GBO1;
wire R18C37_GB70;
wire R28C16_B2;
wire R28C34_E22;
wire R10C34_X01;
wire R9C19_GBO0;
wire R27C24_GB60;
wire R16C20_GT00;
wire R10C19_N80;
wire R3C30_GBO1;
wire R9C42_GT10;
wire R6C37_GBO0;
wire R15C36_GB10;
wire R14C5_GB50;
wire R28C4_B3;
wire R3C21_GB50;
wire R26C29_GT00;
wire R4C44_GB60;
wire R10C26_B4;
wire R4C8_GB10;
wire R23C26_GB70;
wire R28C40_Q5;
wire R5C10_GB70;
wire R1C32_W20;
wire R18C4_GB30;
wire R24C29_GBO1;
wire R5C11_GBO0;
wire R10C19_Q7;
wire R28C25_S83;
wire R26C15_GT00;
wire R28C46_N83;
wire R2C1_GT00;
wire R9C9_GB20;
wire R7C22_GBO0;
wire R8C10_GB20;
wire R7C30_GB00;
wire R21C25_GBO0;
wire R5C43_GB20;
wire R10C31_D2;
wire R10C34_D5;
wire R6C5_GB70;
wire R28C10_LSR1;
wire R26C42_GB20;
wire R6C23_GB40;
wire R15C17_GB70;
wire R6C44_GB50;
wire R22C26_GT00;
wire R28C22_E22;
wire R3C25_GB10;
wire R8C37_GB30;
wire R22C15_GT10;
wire R10C16_F3;
wire R10C26_N26;
wire R29C28_C4;
wire R16C32_GT10;
wire R27C26_GBO1;
wire R7C46_GBO0;
wire R7C38_GB70;
wire R10C27_E22;
wire R8C6_GT10;
wire R24C41_GBO1;
wire R28C10_S10;
wire R17C11_GB70;
wire R5C30_GB00;
wire R21C30_GB10;
wire R27C14_GT00;
wire R14C46_GB60;
wire R20C7_GB70;
wire R10C19_N26;
wire R10C7_SEL0;
wire R3C11_GB60;
wire R11C45_GB60;
wire R28C13_S24;
wire R16C15_GB50;
wire R17C11_GB10;
wire R21C27_GBO0;
wire R28C46_C3;
wire R25C16_GB10;
wire R26C40_GB20;
wire R8C44_GB10;
wire R28C43_SEL0;
wire R26C34_GB20;
wire R25C12_GB60;
wire R22C19_GB50;
wire R13C40_GBO1;
wire R3C33_GB70;
wire R20C8_GBO1;
wire R29C28_E25;
wire R9C28_GB30;
wire R14C33_GB40;
wire R28C22_C6;
wire R7C3_GB50;
wire R11C13_GB40;
wire R20C30_GB60;
wire R10C27_A2;
wire R10C22_N80;
wire R20C7_GB20;
wire R13C8_GT10;
wire R21C6_GBO1;
wire R15C33_GB40;
wire R26C12_GB70;
wire R28C31_N24;
wire R25C27_GB00;
wire R23C33_GB50;
wire R10C37_N24;
wire R16C15_GB10;
wire R4C4_GB50;
wire R23C18_GB10;
wire R1C1_W21;
wire R27C37_GB40;
wire R22C41_GBO0;
wire R10C43_A7;
wire R10C34_N26;
wire R24C30_GB30;
wire R1C47_S27;
wire R29C28_B0;
wire R27C17_GT00;
wire R27C31_GB30;
wire R28C40_W26;
wire R23C11_GBO0;
wire R11C35_GB00;
wire R17C1_GBO1;
wire R7C32_GB50;
wire R17C21_GT00;
wire R10C25_E10;
wire R28C34_N26;
wire R28C28_SEL0;
wire R17C46_GB20;
wire R28C13_D2;
wire R15C10_GT10;
wire R14C45_GT10;
wire R17C46_GB10;
wire R11C37_GBO0;
wire R10C10_W25;
wire R10C37_LSR0;
wire R28C43_E25;
wire R2C29_GBO1;
wire R10C19_D5;
wire R2C36_SPINE4;
wire R10C31_S82;
wire R10C7_X01;
wire R15C39_GT10;
wire R20C22_GB00;
wire R16C21_GT10;
wire R16C39_GB70;
wire R10C7_N11;
wire R12C9_GT00;
wire R28C7_Q5;
wire R23C33_GB30;
wire R24C10_GB30;
wire R23C5_GB20;
wire R24C7_GB60;
wire R20C25_GB40;
wire R27C18_GB20;
wire R18C30_GBO1;
wire R11C38_GB70;
wire R10C26_E26;
wire R10C40_B7;
wire R23C18_GB20;
wire R18C24_GB30;
wire R12C31_GT10;
wire R25C35_GB70;
wire R9C9_GBO1;
wire R26C27_GB10;
wire R27C17_GB30;
wire R8C12_GB50;
wire R4C38_GB50;
wire R15C32_GB40;
wire R28C34_F5;
wire R27C8_GT10;
wire R28C10_N81;
wire R17C11_GB40;
wire R2C39_SPINE1;
wire R9C6_GBO1;
wire R17C28_GB20;
wire R11C23_GB40;
wire R16C3_GBO1;
wire R10C7_C2;
wire R8C34_GBO1;
wire R10C31_Q5;
wire R27C18_GB50;
wire R10C30_B4;
wire R25C41_GT00;
wire R15C8_GB10;
wire R12C18_GB10;
wire R23C46_GB70;
wire R14C42_GB70;
wire R21C8_GB20;
wire R17C24_GB40;
wire R28C13_B3;
wire R10C13_E10;
wire R12C26_GB10;
wire R9C20_GT00;
wire R28C13_N10;
wire R10C16_Q5;
wire R8C37_GB50;
wire R28C43_W12;
wire R18C17_GB60;
wire R2C2_GB20;
wire R18C5_GB10;
wire R10C13_A5;
wire R12C17_GT00;
wire R12C5_GB70;
wire R28C46_A2;
wire R14C14_GB40;
wire R15C32_GB10;
wire R3C22_GBO0;
wire R10C22_W27;
wire R10C37_X04;
wire R16C31_GB50;
wire R12C43_GB50;
wire R2C40_GT00;
wire R11C9_GT00;
wire R14C29_GBO0;
wire R10C43_E13;
wire R11C18_GB00;
wire R12C45_GBO0;
wire R26C36_GB00;
wire R21C5_GBO1;
wire R8C25_GT10;
wire R25C14_GT00;
wire R9C28_GB40;
wire R28C19_E25;
wire R16C46_GB60;
wire R20C35_GB40;
wire R28C28_B0;
wire R9C27_GB60;
wire R20C11_GBO0;
wire R2C7_GT10;
wire R4C34_GT10;
wire R3C4_GB60;
wire R3C44_GB30;
wire R6C25_GT10;
wire R12C15_GT10;
wire R18C6_GB70;
wire R16C34_GB30;
wire R24C26_GBO0;
wire R11C34_GBO1;
wire R27C41_GB70;
wire R10C28_E11;
wire R10C26_D7;
wire R14C30_GB10;
wire R5C41_GB10;
wire R25C19_GBO1;
wire R23C44_GB10;
wire R28C28_CLK0;
wire R14C41_GBO0;
wire R10C25_C3;
wire R21C18_GT00;
wire R18C40_GB60;
wire R28C4_SEL6;
wire R10C16_N80;
wire R28C28_W10;
wire R28C31_B1;
wire R7C28_GB00;
wire R26C35_GB10;
wire R16C37_GBO0;
wire R6C11_GT00;
wire R16C28_GT00;
wire R10C40_S12;
wire R10C27_F5;
wire R22C15_GB30;
wire R4C27_GB40;
wire R14C45_GB20;
wire R20C2_GB10;
wire R20C34_GBO0;
wire R20C2_GB30;
wire R23C7_GB60;
wire R28C7_Q0;
wire R10C27_W20;
wire R28C19_N80;
wire R2C15_GT10;
wire R24C21_GBO1;
wire R10C40_C2;
wire R3C45_GB60;
wire R20C44_GB20;
wire R23C35_GT10;
wire R8C36_GB20;
wire R12C46_GB50;
wire R10C31_W12;
wire R28C34_A2;
wire R2C29_GB20;
wire R18C3_GB30;
wire R28C37_A0;
wire R21C33_GB60;
wire R3C16_GB70;
wire R20C27_GBO0;
wire R18C19_GT00;
wire R13C45_GT10;
wire R21C20_GB50;
wire R15C34_GB30;
wire R28C22_X04;
wire R5C8_GB20;
wire R20C18_GT10;
wire R24C33_GT00;
wire R10C19_CE1;
wire R27C26_GB40;
wire R10C40_X01;
wire R28C46_W21;
wire R10C27_UNK125;
wire R1C1_Q5;
wire R10C29_N82;
wire R27C13_GT10;
wire R7C19_GBO0;
wire R7C2_GBO1;
wire R24C15_GB40;
wire R10C13_S13;
wire R16C33_GBO1;
wire R27C38_GB10;
wire R28C10_N13;
wire R20C10_GB20;
wire R28C46_CE0;
wire R11C14_GB30;
wire R22C43_GB60;
wire R28C19_X05;
wire R21C37_GB40;
wire R9C11_GB40;
wire R28C25_C7;
wire R10C29_B0;
wire R22C36_GB50;
wire R28C34_C2;
wire R10C7_EW10;
wire R17C39_GT10;
wire R27C23_GB40;
wire R14C23_GBO1;
wire R28C16_D4;
wire R11C26_GB40;
wire R10C30_Q0;
wire R18C18_GT10;
wire R9C18_GB60;
wire R23C7_GB10;
wire R4C30_GB50;
wire R26C41_GB70;
wire R12C16_GT10;
wire R9C25_GB00;
wire R28C16_N24;
wire R11C2_GT10;
wire R4C46_GB00;
wire R9C43_GB60;
wire R17C12_GBO1;
wire R11C22_GT00;
wire R10C31_C7;
wire R11C35_GB20;
wire R24C38_GB40;
wire R28C46_SN10;
wire R7C20_GB30;
wire R28C13_S27;
wire R29C28_W25;
wire R23C26_GB10;
wire R8C40_GB40;
wire R21C8_GBO1;
wire R3C44_GBO0;
wire R22C36_GT00;
wire R10C31_N24;
wire R28C37_X08;
wire R29C28_LSR2;
wire R13C21_GB30;
wire R8C5_GBO1;
wire R3C41_GT00;
wire R8C16_GB30;
wire R18C46_GB10;
wire R16C8_GB60;
wire R26C31_GB20;
wire R21C10_GT00;
wire R25C41_GT10;
wire R7C2_GB20;
wire R3C26_GB40;
wire R10C26_E23;
wire R26C42_GT10;
wire R27C45_GB50;
wire R28C19_SEL6;
wire R8C5_GT10;
wire R9C24_GT00;
wire R11C40_GB50;
wire R28C16_SEL7;
wire R22C37_GT10;
wire R28C28_X07;
wire R12C32_GB40;
wire R6C36_GB20;
wire R17C14_GBO1;
wire R15C23_GB30;
wire R4C1_GT10;
wire R13C20_GB20;
wire R23C7_GB30;
wire R4C3_GB60;
wire R24C31_GB10;
wire R8C5_GB70;
wire R13C24_GB10;
wire R21C12_GBO0;
wire R25C9_GB40;
wire R21C17_GBO1;
wire R3C27_GB70;
wire R26C2_GB60;
wire R12C20_GB20;
wire R27C45_GB30;
wire R2C42_GB00;
wire R8C14_GB20;
wire R11C11_GB50;
wire R5C32_GB10;
wire R10C43_W80;
wire R23C32_GB50;
wire R16C9_GT10;
wire R21C20_GB70;
wire R28C19_A3;
wire R14C5_GB70;
wire R9C10_GB60;
wire R13C35_GB10;
wire R26C42_GB70;
wire R14C42_GBO0;
wire R24C45_GB10;
wire R7C10_GB60;
wire R7C22_GB00;
wire R9C21_GB40;
wire R27C10_GB30;
wire R28C40_SEL4;
wire R12C6_GBO1;
wire R28C40_X05;
wire R10C28_Q0;
wire R28C46_C5;
wire R20C38_GB20;
wire R3C15_GB20;
wire R18C17_GT10;
wire R8C20_GB00;
wire R13C16_GB60;
wire R7C34_GB50;
wire R21C14_GB40;
wire R22C16_GBO0;
wire R8C34_GB40;
wire R21C4_GB40;
wire R15C41_GB30;
wire R10C13_N11;
wire R28C13_A6;
wire R10C13_B5;
wire R12C44_GB50;
wire R13C46_GB50;
wire R28C13_N25;
wire R11C9_GB60;
wire R26C39_GB70;
wire R15C23_GB50;
wire R7C39_GB10;
wire R28C16_X05;
wire R11C14_GB10;
wire R11C17_GB10;
wire R9C8_GB00;
wire R2C11_GT00;
wire R26C12_GBO0;
wire R22C40_GT00;
wire R20C39_SPINE29;
wire R28C22_N23;
wire R23C15_GT00;
wire R18C15_GT10;
wire R17C41_GB60;
wire R10C22_F6;
wire R15C42_GB20;
wire R7C28_GB10;
wire R22C24_GB00;
wire R10C19_X01;
wire R28C37_N81;
wire R21C18_GT10;
wire R10C34_E11;
wire R15C41_GB40;
wire R23C11_GB70;
wire R10C34_SEL7;
wire R17C30_GT10;
wire R10C22_S10;
wire R2C45_GB40;
wire R28C16_Q0;
wire R23C23_GB50;
wire R20C2_GT00;
wire R27C14_GB00;
wire R21C12_GBO1;
wire R10C31_F1;
wire R10C40_F3;
wire R1C47_F6;
wire R26C26_GB50;
wire R28C28_E23;
wire R21C45_GB40;
wire R24C36_GB70;
wire R28C25_S23;
wire R1C32_S27;
wire R9C41_GT00;
wire R8C3_GB70;
wire R16C2_GBO1;
wire R3C41_GB20;
wire R26C46_GBO1;
wire R23C14_GB60;
wire R10C25_N13;
wire R14C12_GB50;
wire R13C30_GB40;
wire R13C10_GB00;
wire R10C43_B7;
wire R7C10_GB70;
wire R25C31_GB20;
wire R29C28_SEL4;
wire R3C4_GB50;
wire R11C43_GB00;
wire R10C28_X07;
wire R10C37_S24;
wire R28C19_W13;
wire R7C7_GB60;
wire R8C24_GB50;
wire R25C23_GB00;
wire R11C42_GB60;
wire R10C37_N23;
wire R3C38_GBO0;
wire R18C10_GBO0;
wire R23C42_GB20;
wire R21C34_GB20;
wire R10C16_S81;
wire R28C19_S80;
wire R6C46_GB10;
wire R10C19_SEL3;
wire R16C36_GT00;
wire R28C4_E13;
wire R18C39_GT10;
wire R25C6_GB30;
wire R10C19_C5;
wire R24C23_GB00;
wire R10C34_E23;
wire R6C35_GBO0;
wire R26C42_GB00;
wire R10C22_X02;
wire R6C33_GB10;
wire R5C43_GB50;
wire R10C10_E13;
wire R7C37_GB20;
wire R25C45_GB70;
wire R2C23_GB60;
wire R1C32_C4;
wire R2C7_GB50;
wire R15C10_GB60;
wire R5C37_GBO0;
wire R28C7_SEL7;
wire R20C5_GB70;
wire R18C33_GB20;
wire R9C26_GB20;
wire R1C1_SEL5;
wire R10C27_SPINE8;
wire R5C31_GB70;
wire R4C34_GBO1;
wire R10C7_N20;
wire R10C19_F3;
wire R28C43_C4;
wire R6C4_GT00;
wire R10C43_D7;
wire R2C31_GB20;
wire R10C13_F0;
wire R21C17_GB20;
wire R24C34_GT00;
wire R11C17_GB40;
wire R26C25_GB20;
wire R27C34_GB10;
wire R3C22_GB40;
wire R28C31_N20;
wire R10C7_D3;
wire R21C25_GT00;
wire R26C3_GB70;
wire R3C34_GB70;
wire R5C2_GB10;
wire R5C22_GB70;
wire R14C38_GB60;
wire R4C25_GB40;
wire R22C25_GB00;
wire R15C11_GB50;
wire R25C36_GB20;
wire R10C43_SEL1;
wire R28C4_S22;
wire R26C28_GB60;
wire R3C45_GB70;
wire R23C9_GBO1;
wire R24C13_GB10;
wire R1C32_E83;
wire R17C8_GT10;
wire R1C47_N10;
wire R13C29_GB20;
wire R21C25_GT10;
wire R2C33_GB10;
wire R10C26_Q3;
wire R20C17_GB00;
wire R28C13_Q0;
wire R28C16_N23;
wire R1C47_S25;
wire R28C19_E10;
wire R16C8_GB70;
wire R5C6_GBO1;
wire R12C43_GBO1;
wire R3C12_GT10;
wire R22C8_GB10;
wire R27C30_GB20;
wire R16C35_GB30;
wire R15C28_GT00;
wire R13C12_GB20;
wire R25C19_GB70;
wire R10C19_LSR1;
wire R14C32_GT00;
wire R20C10_GB10;
wire R3C5_GT00;
wire R18C35_GB70;
wire R10C13_D1;
wire R26C10_GB70;
wire R22C26_GT10;
wire R24C33_GB70;
wire R9C26_GB50;
wire R8C36_GB60;
wire R28C10_X01;
wire R21C37_GB60;
wire R27C6_GT10;
wire R22C30_GB40;
wire R28C31_E25;
wire R15C4_GT00;
wire R4C35_GBO0;
wire R21C45_GT10;
wire R3C11_GT10;
wire R17C28_GB70;
wire R14C7_GB10;
wire R28C16_E10;
wire R28C19_F5;
wire R5C1_GT00;
wire R10C10_N82;
wire R28C4_D6;
wire R27C40_GB70;
wire R28C13_C2;
wire R14C39_GB40;
wire R20C33_GT00;
wire R3C10_GB20;
wire R9C29_GB40;
wire R25C6_GBO1;
wire R15C25_GB30;
wire R10C26_LSR0;
wire R10C40_N80;
wire R11C5_GT10;
wire R11C37_GB60;
wire R2C30_SPINE2;
wire R17C31_GT00;
wire R14C20_GB40;
wire R4C40_GB50;
wire R6C34_GB70;
wire R14C30_GB20;
wire R16C24_GB40;
wire R24C39_GB60;
wire R5C5_GB10;
wire R28C40_E24;
wire R10C10_SEL0;
wire R22C6_GT10;
wire R10C22_B6;
wire R28C25_A1;
wire R22C25_GT10;
wire R12C26_GB20;
wire R3C31_GBO1;
wire R10C43_W82;
wire R10C13_LSR0;
wire R10C27_E83;
wire R20C3_GT10;
wire R10C7_W10;
wire R28C7_SEL2;
wire R20C24_SPINE20;
wire R9C27_GBO1;
wire R12C8_GB40;
wire R28C25_E25;
wire R7C32_GT00;
wire R5C33_GB00;
wire R10C37_E26;
wire R28C13_CLK2;
wire R24C17_GT10;
wire R27C26_GT00;
wire R18C15_GB40;
wire R24C4_GB50;
wire R28C43_W81;
wire R12C22_GBO0;
wire R14C18_GB20;
wire R11C22_GB30;
wire R4C28_GB00;
wire R7C25_GT00;
wire R18C1_GT00;
wire R24C45_GT10;
wire R26C22_GBO0;
wire R24C27_GB70;
wire R1C28_CLK0;
wire R10C22_W25;
wire R6C9_GB50;
wire R28C28_X04;
wire R28C7_D2;
wire R28C10_CE2;
wire R26C46_GB70;
wire R12C41_GB70;
wire R10C30_A0;
wire R13C21_GT10;
wire R14C42_GB40;
wire R12C10_GB40;
wire R20C32_GB00;
wire R6C38_GB70;
wire R10C19_S23;
wire R10C16_B3;
wire R23C31_GB40;
wire R17C3_GB20;
wire R17C27_GT00;
wire R5C29_GBO1;
wire R24C21_GB50;
wire R10C25_A2;
wire R10C29_N12;
wire R17C41_GT10;
wire R28C43_E83;
wire R18C5_GB00;
wire R13C13_GBO0;
wire R8C13_GB20;
wire R5C9_GB40;
wire R17C24_GB20;
wire R20C12_GB70;
wire R9C31_GB50;
wire R23C39_GBO1;
wire R28C13_N20;
wire R28C13_D7;
wire R10C30_UNK124;
wire R8C41_GT00;
wire R5C10_GB00;
wire R14C10_GB60;
wire R20C34_GB40;
wire R28C46_B4;
wire R21C29_GB00;
wire R21C43_GB00;
wire R12C40_GB30;
wire R10C25_N83;
wire R11C37_GB40;
wire R15C37_GB30;
wire R18C3_GT10;
wire R21C29_GB30;
wire R23C43_GBO1;
wire R28C34_N10;
wire R28C28_S20;
wire R3C13_GBO0;
wire R6C42_GB00;
wire R28C37_X07;
wire R18C7_GB40;
wire R27C46_GT00;
wire R20C16_SPINE16;
wire R11C18_GT10;
wire R8C1_GT10;
wire R6C15_GBO1;
wire R10C31_N13;
wire R4C11_GT00;
wire R28C13_SN10;
wire R28C28_F7;
wire R20C30_GT10;
wire R23C15_GB50;
wire R24C23_GB40;
wire R23C9_GB70;
wire R28C46_N12;
wire R10C28_W20;
wire R28C40_E22;
wire R6C38_GT00;
wire R3C38_GB30;
wire R24C16_GB70;
wire R24C19_GT00;
wire R13C30_GB00;
wire R24C5_GT00;
wire R28C28_Q6;
wire R16C35_GBO1;
wire R9C38_GT10;
wire R21C18_GB70;
wire R10C29_EW20;
wire R10C43_X08;
wire R4C6_GB70;
wire R9C33_GT10;
wire R20C15_GT00;
wire R9C20_GB70;
wire R13C5_GB10;
wire R3C40_GB70;
wire R27C34_GBO1;
wire R20C43_GB70;
wire R10C31_B4;
wire R12C5_GBO1;
wire R26C44_GB60;
wire R14C39_GBO0;
wire R1C47_W21;
wire R8C11_GBO0;
wire R13C42_GT10;
wire R7C18_GB00;
wire R25C40_GB00;
wire R11C27_GB10;
wire R28C34_F7;
wire R10C31_E27;
wire R28C16_S13;
wire R28C43_C6;
wire R7C3_GT00;
wire R27C6_GB30;
wire R15C11_GB30;
wire R23C4_GB20;
wire R22C27_GB30;
wire R21C7_GB40;
wire R12C28_GB30;
wire R16C19_GB70;
wire R6C45_GB50;
wire R5C17_GB10;
wire R4C25_GB70;
wire R26C17_GB70;
wire R16C39_GB40;
wire R10C19_N25;
wire R10C29_CE1;
wire R28C46_Q1;
wire R10C10_S24;
wire R10C27_S24;
wire R28C37_B4;
wire R13C29_GB50;
wire R24C11_GB40;
wire R10C43_N26;
wire R28C4_A6;
wire R28C10_A0;
wire R25C27_GT10;
wire R28C31_N83;
wire R28C13_C0;
wire R16C32_GB70;
wire R15C15_GB60;
wire R22C37_GB70;
wire R3C15_GB00;
wire R2C45_GB30;
wire R23C36_GT10;
wire R12C45_GB50;
wire R20C7_SPINE17;
wire R13C45_GBO0;
wire R25C2_GB70;
wire R11C42_GB00;
wire R17C37_GT10;
wire R3C1_GT00;
wire R10C29_A4;
wire R22C17_GB30;
wire R12C46_GT10;
wire R28C16_F6;
wire R9C7_GB00;
wire R28C13_E22;
wire R22C4_GB70;
wire R7C11_GBO1;
wire R5C4_GT00;
wire R18C46_GT10;
wire R3C30_GB20;
wire R15C37_GB10;
wire R9C39_GT00;
wire R27C33_GB20;
wire R22C20_GB30;
wire R4C43_GT10;
wire R1C47_C1;
wire R29C28_Q6;
wire R26C2_GB30;
wire R12C3_GB60;
wire R28C13_D4;
wire R14C40_GT00;
wire R7C21_GB60;
wire R24C41_GB60;
wire R14C3_GB50;
wire R27C33_GBO1;
wire R6C38_GB30;
wire R3C8_GBO1;
wire R4C43_GB40;
wire R10C16_A5;
wire R13C7_GT10;
wire R2C15_GB60;
wire R28C46_X02;
wire R10C7_SEL1;
wire R26C18_GB10;
wire R14C15_GB30;
wire R10C13_S22;
wire R20C43_GB40;
wire R28C34_X01;
wire R3C24_GB70;
wire R11C33_GB40;
wire R15C23_GB20;
wire R1C32_S82;
wire R5C39_GB50;
wire R10C40_E26;
wire R10C29_UNK123;
wire R26C43_GB30;
wire R13C19_GB00;
wire R10C30_CLK2;
wire R28C4_W10;
wire R27C14_GBO1;
wire R11C4_GB40;
wire R28C25_N22;
wire R10C40_F0;
wire R21C33_GB50;
wire R10C37_SEL4;
wire R14C11_GB10;
wire R26C12_GB00;
wire R17C37_GB50;
wire R23C42_GB50;
wire R10C7_LSR0;
wire R1C28_SEL1;
wire R8C31_GB20;
wire R3C34_GB10;
wire R15C36_GB00;
wire R6C6_GB30;
wire R8C44_GT10;
wire R25C25_GB00;
wire R23C22_GB20;
wire R25C45_GB20;
wire R10C40_EW20;
wire R10C26_CE2;
wire R11C4_GT10;
wire R9C42_GB00;
wire R14C43_GT00;
wire R4C15_GB60;
wire R26C37_GT00;
wire R5C22_GBO0;
wire R2C23_GB30;
wire R18C28_GB40;
wire R7C31_GT10;
wire R5C37_GB30;
wire R9C40_GB00;
wire R28C40_N12;
wire R24C11_GT10;
wire R2C22_GBO0;
wire R21C44_GBO1;
wire R7C28_GT10;
wire R17C6_GB00;
wire R27C20_GB10;
wire R20C1_GBO0;
wire R13C12_GB60;
wire R3C42_GB30;
wire R10C28_UNK122;
wire R27C33_GB60;
wire R24C20_GB00;
wire R5C2_GBO1;
wire R14C36_GT10;
wire R28C7_N20;
wire R5C33_GB60;
wire R21C45_GB20;
wire R25C33_GB00;
wire R23C43_GB10;
wire R25C22_GB20;
wire R6C14_GBO0;
wire R18C38_GB60;
wire R1C1_D1;
wire R13C11_GT00;
wire R7C42_GBO1;
wire R12C33_GBO0;
wire R3C29_GB40;
wire R20C16_GT00;
wire R29C28_X01;
wire R5C43_GT10;
wire R22C12_GB00;
wire R13C41_GB30;
wire R10C31_W80;
wire R5C32_GB60;
wire R6C18_GB70;
wire R23C22_GB40;
wire R28C22_W81;
wire R6C10_GB50;
wire R10C16_S20;
wire R4C13_GB40;
wire R20C7_GB30;
wire R28C40_SEL5;
wire R15C34_GB50;
wire R6C32_GB20;
wire R5C38_GBO1;
wire R1C1_E11;
wire R24C30_GB60;
wire R13C42_GB10;
wire R9C2_GB70;
wire R2C9_GT10;
wire R11C27_GT10;
wire R10C25_LSR0;
wire R21C35_GBO0;
wire R20C8_GB70;
wire R8C42_GBO0;
wire R10C22_C1;
wire R20C19_GB60;
wire R2C31_GB50;
wire R27C41_GBO0;
wire R14C4_GB00;
wire R11C14_GT10;
wire R21C42_GB10;
wire R17C29_GB30;
wire R27C43_GB30;
wire R1C47_D7;
wire R28C37_C7;
wire R28C28_N13;
wire R28C46_LSR1;
wire R24C19_GB50;
wire R20C1_SPINE19;
wire R25C29_GT10;
wire R4C35_GB60;
wire R9C13_GB10;
wire R7C6_GB10;
wire R12C16_GB10;
wire R10C43_F4;
wire R2C20_GB20;
wire R23C19_GBO1;
wire R8C19_GT00;
wire R6C29_GBO1;
wire R20C36_GBO0;
wire R10C16_LSR2;
wire R5C33_GBO1;
wire R1C1_E27;
wire R9C13_GBO0;
wire R6C5_GB00;
wire R14C32_GB60;
wire R10C34_E22;
wire R8C18_GBO0;
wire R24C8_GB70;
wire R9C8_GB20;
wire R23C21_GB70;
wire R23C26_GB40;
wire R20C41_GB00;
wire R5C5_GT10;
wire R12C25_GB70;
wire R24C36_GB10;
wire R10C34_F2;
wire R24C8_GT10;
wire R28C28_E26;
wire R28C40_E12;
wire R10C28_E81;
wire R28C37_S82;
wire R6C3_GT00;
wire R28C37_N11;
wire R5C30_GB10;
wire R10C13_CE2;
wire R28C31_S10;
wire R24C30_GT10;
wire R14C44_GT10;
wire R3C28_GB60;
wire R9C23_GT00;
wire R7C27_GT10;
wire R22C9_GB70;
wire R14C44_GB10;
wire R28C28_W11;
wire R28C34_SEL2;
wire R12C20_GT10;
wire R11C41_GB60;
wire R9C5_GB60;
wire R18C25_GBO1;
wire R6C42_GB10;
wire R2C6_GB20;
wire R10C30_B6;
wire R2C27_GB00;
wire R7C7_GT10;
wire R26C29_GB00;
wire R10C7_W21;
wire R13C19_GB10;
wire R10C40_CE2;
wire R24C7_GB00;
wire R22C2_GB10;
wire R4C4_GB10;
wire R13C23_GB70;
wire R13C24_GT10;
wire R20C23_GBO1;
wire R22C41_GBO1;
wire R5C23_GB00;
wire R7C24_GB20;
wire R10C28_A7;
wire R18C16_GBO0;
wire R11C26_GB00;
wire R23C36_GB40;
wire R1C1_X05;
wire R10C7_D5;
wire R28C13_E23;
wire R17C26_GB50;
wire R12C39_GT10;
wire R12C14_GB20;
wire R8C4_GB30;
wire R17C9_GB20;
wire R29C28_E81;
wire R10C29_S80;
wire R14C13_GB60;
wire R16C41_GB10;
wire R28C31_SEL7;
wire R5C28_GB40;
wire R28C19_A6;
wire R6C7_GB20;
wire R28C43_E11;
wire R12C21_GT10;
wire R28C13_N12;
wire R8C13_GT00;
wire R28C25_S13;
wire R12C33_GT10;
wire R10C19_B4;
wire R5C32_GB20;
wire R10C19_X07;
wire R4C1_GBO0;
wire R1C47_N27;
wire R14C45_GB50;
wire R11C8_GB70;
wire R28C34_A5;
wire R28C19_SEL2;
wire R26C34_GT10;
wire R11C27_GB60;
wire R18C13_GB00;
wire R7C39_GB60;
wire R25C20_GB10;
wire R16C27_GB10;
wire R2C14_SPINE10;
wire R28C13_E81;
wire R4C14_GB70;
wire R2C45_GB00;
wire R13C27_GBO0;
wire R10C26_SEL2;
wire R10C27_N13;
wire R8C25_GB60;
wire R16C8_GB30;
wire R25C27_GB40;
wire R25C36_GB60;
wire R4C20_GB20;
wire R27C21_GT10;
wire R24C5_GBO1;
wire R28C16_E27;
wire R5C28_GB50;
wire R8C22_GB70;
wire R6C8_GB40;
wire R2C43_GT10;
wire R15C33_GT10;
wire R5C9_GB00;
wire R1C28_F6;
wire R25C19_GB60;
wire R16C7_GT10;
wire R15C26_GB40;
wire R21C33_GB30;
wire R12C12_GB20;
wire R11C37_GB30;
wire R27C35_GB00;
wire R23C34_GB40;
wire R28C19_D2;
wire R25C44_GB40;
wire R26C46_GBO0;
wire R28C34_S80;
wire R10C40_W10;
wire R10C10_N12;
wire R28C43_S24;
wire R28C19_Q6;
wire R10C28_F7;
wire R5C12_GT00;
wire R2C34_GT10;
wire R12C4_GBO1;
wire R3C33_GT10;
wire R17C23_GBO0;
wire R27C29_GB50;
wire R2C22_GB40;
wire R22C6_GB70;
wire R28C10_A2;
wire R11C14_GBO1;
wire R3C46_GB60;
wire R11C4_GB30;
wire R6C11_GB60;
wire R5C17_GB60;
wire R6C41_GT00;
wire R25C41_GB00;
wire R12C13_GB20;
wire R3C17_GB40;
wire R10C34_S83;
wire R10C34_S12;
wire R13C15_GB10;
wire R16C29_GB20;
wire R6C3_GB20;
wire R27C44_GB20;
wire R15C3_GBO1;
wire R22C24_GB40;
wire R12C9_GBO0;
wire R13C20_GT00;
wire R28C40_S11;
wire R20C10_GB50;
wire R3C4_GB40;
wire R8C8_GB20;
wire R28C13_CE1;
wire R7C7_GB70;
wire R10C40_C3;
wire R5C40_GB10;
wire R28C31_B2;
wire R27C27_GB60;
wire R25C8_GB70;
wire R25C19_GB50;
wire R20C37_GB10;
wire R10C37_W27;
wire R28C43_S21;
wire R13C10_GB60;
wire R18C20_GBO0;
wire R9C30_GB20;
wire R10C7_S80;
wire R5C27_GT10;
wire R28C22_A7;
wire R25C36_GB30;
wire R22C29_GBO1;
wire R14C38_GB10;
wire R14C9_GT00;
wire R17C12_GB10;
wire R24C41_GT00;
wire R18C38_GB30;
wire R16C42_GBO1;
wire R5C6_GT00;
wire R10C13_W81;
wire R24C19_GB10;
wire R18C40_GB30;
wire R5C46_GB70;
wire R20C39_GB40;
wire R2C22_GB70;
wire R18C29_GB40;
wire R21C5_GB10;
wire R5C35_GBO1;
wire R28C4_SEL1;
wire R25C3_GT10;
wire R12C32_GB70;
wire R28C4_CE2;
wire R10C7_S23;
wire R17C6_GT10;
wire R10C7_Q2;
wire R13C44_GB10;
wire R10C34_A4;
wire R25C29_GB00;
wire R10C10_A1;
wire R9C44_GT00;
wire R10C13_X06;
wire R8C25_GB00;
wire R1C28_CLK1;
wire R23C15_GB00;
wire R18C18_GB30;
wire R17C29_GB70;
wire R27C20_GBO0;
wire R16C40_GB60;
wire R8C31_GB60;
wire R7C12_GBO1;
wire R24C46_GB40;
wire R11C23_GT10;
wire R5C12_GB10;
wire R2C45_SPINE3;
wire R26C4_GBO0;
wire R27C24_GB70;
wire R12C30_GT10;
wire R25C27_GB30;
wire R16C42_GBO0;
wire R1C47_A3;
wire R4C42_GB60;
wire R10C31_W82;
wire R7C43_GB20;
wire R20C41_GB20;
wire R10C19_A7;
wire R9C10_GB40;
wire R15C20_GBO0;
wire R10C19_F0;
wire R9C14_GBO0;
wire R28C43_F0;
wire R23C9_GT10;
wire R15C9_GB10;
wire R3C31_GB10;
wire R21C2_GT00;
wire R18C27_GBO0;
wire R28C7_W22;
wire R9C44_GBO1;
wire R22C16_GB70;
wire R10C28_Q6;
wire R24C40_GB30;
wire R15C24_GBO1;
wire R10C28_E10;
wire R15C43_GT00;
wire R17C15_GB10;
wire R20C23_GB50;
wire R18C7_GB10;
wire R1C32_Q3;
wire R27C19_GB10;
wire R14C21_GB30;
wire R10C31_Q2;
wire R12C43_GT00;
wire R28C43_C7;
wire R6C21_GB50;
wire R15C18_GT10;
wire R5C34_GB50;
wire R17C27_GBO0;
wire R10C22_S11;
wire R2C14_GB10;
wire R12C7_GB10;
wire R9C16_GB50;
wire R25C14_GB00;
wire R3C25_GB00;
wire R24C40_GBO0;
wire R21C26_GT00;
wire R16C12_GB50;
wire R7C31_GB00;
wire R23C14_GBO1;
wire R3C6_GB10;
wire R27C7_GB70;
wire R20C5_GBO0;
wire R10C43_B3;
wire R26C27_GB20;
wire R8C38_GB70;
wire R4C46_GB30;
wire R5C25_GB40;
wire R22C12_GT00;
wire R18C36_GB20;
wire R9C8_GB70;
wire R20C11_SPINE17;
wire R5C38_GB00;
wire R28C43_W27;
wire R20C31_SPINE29;
wire R18C41_GB50;
wire R2C2_GB10;
wire R2C22_GB30;
wire R28C31_B4;
wire R27C39_GB50;
wire R22C31_GB10;
wire R8C31_GB40;
wire R28C40_E11;
wire R18C39_GB30;
wire R11C28_GT10;
wire R6C41_GB20;
wire R15C9_GBO1;
wire R28C7_D6;
wire R28C25_W24;
wire R9C28_GB10;
wire R3C11_GB20;
wire R17C10_GB50;
wire R17C5_GB50;
wire R14C29_GB00;
wire R27C42_GB70;
wire R18C28_GB60;
wire R15C26_GBO0;
wire R28C46_S27;
wire R3C37_GB70;
wire R20C23_GB40;
wire R24C43_GB10;
wire R21C36_GT10;
wire R23C29_GB00;
wire R9C15_GBO0;
wire R7C35_GB40;
wire R10C25_Q1;
wire R10C30_SEL3;
wire R8C4_GB20;
wire R1C47_F5;
wire R16C6_GB20;
wire R9C4_GT10;
wire R26C23_GB30;
wire R21C5_GB40;
wire R7C14_GT10;
wire R26C33_GB00;
wire R27C30_GB00;
wire R18C17_GB30;
wire R24C40_GB00;
wire R10C30_E27;
wire R11C46_GB70;
wire R21C10_GB00;
wire R3C32_GB60;
wire R10C22_S81;
wire R10C28_S81;
wire R10C43_Q7;
wire R21C23_GBO1;
wire R23C28_GB70;
wire R10C16_N11;
wire R12C36_GT00;
wire R10C30_D7;
wire R16C13_GB70;
wire R12C18_GT00;
wire R27C10_GBO1;
wire R4C33_GBO0;
wire R14C41_GB10;
wire R28C34_D3;
wire R7C22_GB60;
wire R16C10_GB60;
wire R9C36_GBO0;
wire R25C2_GT00;
wire R27C30_GB50;
wire R15C8_GB00;
wire R10C7_SEL5;
wire R16C17_GB20;
wire R15C14_GB40;
wire R18C7_GT00;
wire R12C41_GT00;
wire R10C26_S10;
wire R2C19_GB60;
wire R17C46_GB50;
wire R10C27_F6;
wire R21C43_GB70;
wire R28C4_E25;
wire R2C2_SPINE10;
wire R10C30_Q1;
wire R24C30_GBO1;
wire R25C18_GB20;
wire R7C2_GB40;
wire R8C40_GBO0;
wire R9C23_GBO0;
wire R18C23_GT00;
wire R17C15_GBO0;
wire R23C25_GB10;
wire R22C12_GB20;
wire R12C17_GB20;
wire R9C30_GB10;
wire R14C4_GT00;
wire R15C29_GB10;
wire R8C42_GB20;
wire R17C19_GB70;
wire R28C28_W21;
wire R24C7_GB30;
wire R27C45_GB00;
wire R23C30_GB10;
wire R21C15_GT00;
wire R11C20_GT00;
wire R28C37_F2;
wire R6C13_GB40;
wire R15C5_GB30;
wire R10C27_LSR2;
wire R4C30_GT00;
wire R16C30_GT00;
wire R13C36_GB70;
wire R10C16_W11;
wire R10C28_X05;
wire R12C24_GT00;
wire R12C14_GT00;
wire R7C43_GB60;
wire R10C16_E22;
wire R24C29_GB20;
wire R25C32_GB70;
wire R2C32_GB00;
wire R26C37_GB40;
wire R6C6_GT10;
wire R10C16_A7;
wire R10C28_D5;
wire R28C16_S25;
wire R12C40_GB00;
wire R9C15_GB40;
wire R13C17_GBO0;
wire R10C37_W21;
wire R23C39_GB60;
wire R21C22_GBO1;
wire R4C44_GB00;
wire R9C39_GB30;
wire R2C17_GB70;
wire R17C38_GB00;
wire R28C31_F1;
wire R29C28_W22;
wire R9C14_GT00;
wire R27C4_GBO1;
wire R24C16_GB20;
wire R11C9_GB40;
wire R11C24_GBO1;
wire R27C31_GB40;
wire R17C31_GB60;
wire R27C8_GT00;
wire R10C34_CE2;
wire R5C22_GT10;
wire R15C28_GB00;
wire R21C9_GB20;
wire R14C9_GB10;
wire R25C8_GT00;
wire R9C1_GT00;
wire R22C14_GBO0;
wire R27C24_GBO1;
wire R28C43_X07;
wire R24C44_GB60;
wire R12C3_GB50;
wire R14C20_GB60;
wire R27C8_GB20;
wire R9C23_GB20;
wire R27C18_GB40;
wire R5C33_GT10;
wire R26C15_GB50;
wire R10C28_SEL5;
wire R10C30_E11;
wire R13C25_GB00;
wire R4C41_GB00;
wire R28C10_EW20;
wire R28C31_E11;
wire R14C25_GBO1;
wire R18C37_GB60;
wire R27C25_GBO1;
wire R2C25_SPINE11;
wire R21C13_GT10;
wire R6C45_GB70;
wire R12C31_GB40;
wire R9C35_GB30;
wire R28C25_SN10;
wire R11C13_GT00;
wire R22C37_GT00;
wire R22C8_GB70;
wire R2C12_GB10;
wire R3C33_GB50;
wire R28C25_SEL1;
wire R27C2_GB70;
wire R12C35_GB20;
wire R28C37_S12;
wire R26C3_GB30;
wire R3C30_GB40;
wire R28C7_S25;
wire R28C43_SEL2;
wire R18C39_GB10;
wire R28C25_N27;
wire R4C45_GB50;
wire R13C8_GB70;
wire R21C32_GB20;
wire R25C23_GBO0;
wire R10C7_A7;
wire R3C12_GB50;
wire R10C7_E26;
wire R16C3_GB70;
wire R9C1_F6;
wire R21C29_GB70;
wire R10C37_E24;
wire R2C43_GB70;
wire R6C23_GBO1;
wire R28C43_W80;
wire R9C3_GB50;
wire R24C18_GB60;
wire R28C34_W81;
wire R3C44_GB10;
wire R10C7_SEL4;
wire R10C27_E80;
wire R28C25_Q3;
wire R10C25_SEL1;
wire R8C14_GT00;
wire R29C28_SEL0;
wire R28C19_F6;
wire R7C34_GB60;
wire R1C1_SN20;
wire R8C4_GB70;
wire R12C35_GB40;
wire R24C40_GB70;
wire R28C7_N80;
wire R24C22_GB10;
wire R15C27_GB20;
wire R14C12_GBO0;
wire R15C6_GT00;
wire R17C37_GB30;
wire R15C41_GT10;
wire R12C18_GB40;
wire R28C25_E13;
wire R23C44_GB40;
wire R7C21_GB40;
wire R10C26_S23;
wire R13C41_GBO1;
wire R28C46_X01;
wire R23C38_GB00;
wire R8C10_GB30;
wire R8C23_GBO1;
wire R4C31_GB30;
wire R13C40_GB10;
wire R29C28_N22;
wire R18C8_GB10;
wire R25C1_GBO0;
wire R17C32_GB20;
wire R10C19_C3;
wire R2C45_GT00;
wire R14C18_GB30;
wire R27C8_GBO1;
wire R23C12_GBO1;
wire R23C41_GB40;
wire R28C19_EW20;
wire R16C45_GB60;
wire R15C3_GT00;
wire R20C9_GB10;
wire R28C10_W20;
wire R8C39_GB10;
wire R10C16_N83;
wire R4C32_GT10;
wire R10C25_X08;
wire R2C30_GT00;
wire R14C31_GB60;
wire R4C24_GB10;
wire R10C29_E23;
wire R20C18_GT00;
wire R3C15_GBO0;
wire R25C32_GB30;
wire R12C34_GB60;
wire R28C13_Q1;
wire R2C27_GB30;
wire R26C23_GT10;
wire R13C14_GT00;
wire R24C43_GB20;
wire R6C18_GBO0;
wire R28C40_E13;
wire R7C35_GB50;
wire R2C5_GT00;
wire R10C30_A4;
wire R15C25_GT00;
wire R4C2_GB00;
wire R7C16_GT10;
wire R29C28_S81;
wire R23C40_GB70;
wire R5C5_GB50;
wire R29C28_E24;
wire R20C19_GT00;
wire R14C19_GB20;
wire R26C34_GB60;
wire R4C34_GB20;
wire R3C18_GT00;
wire R24C7_GB70;
wire R9C45_GB70;
wire R4C7_GB40;
wire R22C41_GB20;
wire R6C10_GB30;
wire R28C7_E24;
wire R4C22_GBO1;
wire R24C10_GB40;
wire R23C39_GB10;
wire R2C15_GBO0;
wire R3C44_GB50;
wire R10C13_E12;
wire R15C23_GB00;
wire R14C13_GB20;
wire R23C3_GB30;
wire R10C27_SPINE9;
wire R27C15_GB10;
wire R20C19_GB70;
wire R7C34_GBO1;
wire R4C22_GT00;
wire R27C4_GBO0;
wire R14C6_GBO0;
wire R28C13_W20;
wire R16C25_GB10;
wire R10C16_N13;
wire R10C16_N25;
wire R26C41_GB60;
wire R28C28_CE1;
wire R11C29_GB30;
wire R25C22_GT10;
wire R28C34_D4;
wire R18C43_GBO1;
wire R16C22_GB70;
wire R10C25_EW20;
wire R17C21_GB30;
wire R2C24_GB30;
wire R13C9_GB60;
wire R2C16_GB40;
wire R7C2_GB10;
wire R10C40_B6;
wire R28C16_EW20;
wire R6C20_GBO1;
wire R18C15_GB10;
wire R15C45_GB00;
wire R21C12_GT00;
wire R12C9_GB40;
wire R1C32_N10;
wire R8C10_GB40;
wire R20C30_GB50;
wire R10C10_D0;
wire R14C10_GB40;
wire R2C25_GB50;
wire R18C29_GT00;
wire R11C40_GBO1;
wire R10C22_W22;
wire R6C20_GB20;
wire R28C37_N27;
wire R20C41_GB40;
wire R5C11_GT10;
wire R17C34_GB10;
wire R12C30_GB30;
wire R26C37_GBO0;
wire R10C10_E25;
wire R16C22_GB30;
wire R21C20_GB00;
wire R8C29_GB60;
wire R27C29_GBO1;
wire R24C42_GT10;
wire R22C24_GB50;
wire R8C33_GB00;
wire R12C13_GB00;
wire R6C32_GBO1;
wire R23C33_GB40;
wire R10C19_S81;
wire R18C24_GBO1;
wire R15C29_GBO1;
wire R13C34_GB10;
wire R28C4_S20;
wire R14C41_GB50;
wire R11C12_GB70;
wire R14C34_GB60;
wire R28C10_D2;
wire R10C40_Q2;
wire R20C4_GBO1;
wire R22C7_GB20;
wire R21C11_GT10;
wire R20C7_GB50;
wire R3C32_GBO0;
wire R1C32_C6;
wire R28C7_D0;
wire R16C22_GBO0;
wire R8C38_GBO1;
wire R4C41_GBO1;
wire R17C2_GB40;
wire R3C18_GB10;
wire R7C16_GB40;
wire R10C28_C6;
wire R17C12_GB40;
wire R21C35_GB20;
wire R17C43_GBO1;
wire R20C28_GB10;
wire R20C10_GB40;
wire R26C40_GT10;
wire R17C45_GBO0;
wire R17C13_GB70;
wire R12C37_GT00;
wire R28C46_SEL2;
wire R28C34_N83;
wire R2C15_GB40;
wire R24C35_GB50;
wire R20C40_GB30;
wire R25C12_GT00;
wire R25C37_GT10;
wire R4C14_GB50;
wire R18C11_GB30;
wire R11C24_GB70;
wire R10C13_N22;
wire R28C4_S25;
wire R28C10_A5;
wire R28C19_N13;
wire R14C29_GB70;
wire R3C35_GT00;
wire R2C12_GB40;
wire R17C18_GB10;
wire R3C44_GBO1;
wire R9C16_GB70;
wire R10C19_F4;
wire R10C28_A1;
wire R5C2_GB00;
wire R11C39_GB30;
wire R28C43_S12;
wire R5C17_GB30;
wire R24C21_GB10;
wire R25C23_GB30;
wire R7C12_GB60;
wire R25C18_GBO1;
wire R25C9_GB60;
wire R8C11_GB20;
wire R22C9_GB00;
wire R25C8_GB00;
wire R26C36_GBO0;
wire R28C22_A4;
wire R14C40_GB60;
wire R28C16_E12;
wire R20C34_GB30;
wire R10C22_N83;
wire R8C21_GB60;
wire R13C19_GB60;
wire R14C35_GB10;
wire R22C7_GB00;
wire R11C10_GB60;
wire R6C14_GT10;
wire R22C38_GB40;
wire R10C30_SPINE5;
wire R7C20_GB70;
wire R2C19_GB20;
wire R20C6_GB60;
wire R7C9_GBO0;
wire R22C15_GB00;
wire R20C38_SPINE26;
wire R22C11_GT10;
wire R27C14_GB70;
wire R2C13_GB30;
wire R7C30_GT00;
wire R13C31_GB00;
wire R16C46_GB00;
wire R20C46_GBO0;
wire R5C5_GBO1;
wire R24C42_GB50;
wire R10C37_E10;
wire R15C44_GBO1;
wire R6C19_GBO0;
wire R15C18_GB40;
wire R2C29_SPINE3;
wire R23C16_GB30;
wire R2C45_GB20;
wire R20C33_GB60;
wire R28C13_E82;
wire R22C40_GB00;
wire R10C10_CLK1;
wire R26C41_GB10;
wire R25C32_GB10;
wire R24C36_GB20;
wire R28C22_SEL4;
wire R2C41_GB50;
wire R15C39_GB60;
wire R3C27_GT10;
wire R9C22_GB70;
wire R28C13_SEL0;
wire R23C18_GB30;
wire R2C3_GBO0;
wire R10C43_E83;
wire R16C22_GB10;
wire R6C46_GB00;
wire R10C13_SEL3;
wire R2C46_GB60;
wire R6C19_GT00;
wire R18C40_GB50;
wire R14C18_GB40;
wire R18C46_GB50;
wire R8C7_GB30;
wire R22C5_GT10;
wire R3C34_GB60;
wire R27C23_GBO0;
wire R13C32_GB10;
wire R27C20_GB40;
wire R10C26_D2;
wire R28C40_X08;
wire R17C38_GT00;
wire R7C19_GT10;
wire R22C4_GB10;
wire R11C8_GB60;
wire R6C44_GB70;
wire R23C46_GB00;
wire R21C43_GBO0;
wire R12C35_GB50;
wire R27C30_GB70;
wire R13C15_GB60;
wire R21C21_GB70;
wire R1C47_B5;
wire R6C19_GB40;
wire R16C30_GB30;
wire R10C7_B0;
wire R11C16_GB00;
wire R5C38_GB50;
wire R3C20_GB10;
wire R8C7_GB60;
wire R28C34_W10;
wire R21C13_GB00;
wire R4C35_GB70;
wire R7C38_GB20;
wire R28C40_B6;
wire R17C28_GB10;
wire R28C4_X07;
wire R9C29_GBO0;
wire R4C39_GB40;
wire R7C18_GB70;
wire R25C39_GB40;
wire R25C37_GB50;
wire R28C37_E82;
wire R20C12_GB50;
wire R6C46_GB20;
wire R27C40_GB30;
wire R6C7_GB40;
wire R3C12_GB00;
wire R17C45_GB70;
wire R7C3_GB10;
wire R10C43_X06;
wire R25C10_GBO1;
wire R25C3_GBO1;
wire R3C25_GB60;
wire R15C21_GBO1;
wire R26C36_GB50;
wire R18C8_GBO0;
wire R11C33_GB10;
wire R4C42_GBO1;
wire R10C22_E10;
wire R10C34_N22;
wire R10C30_E23;
wire R28C7_LSR2;
wire R26C39_GB60;
wire R5C36_GB70;
wire R2C15_GB00;
wire R21C25_GBO1;
wire R9C36_GB60;
wire R10C30_B1;
wire R8C12_GBO1;
wire R27C14_GB40;
wire R15C15_GT00;
wire R21C44_GB30;
wire R23C28_GB60;
wire R13C17_GB70;
wire R24C38_GB20;
wire R10C43_D0;
wire R29C28_B5;
wire R9C34_GB20;
wire R10C37_F4;
wire R18C44_GBO1;
wire R8C13_GBO0;
wire R15C30_GT00;
wire R17C26_GB70;
wire R18C17_GT00;
wire R2C19_SPINE9;
wire R28C46_B6;
wire R3C10_GBO1;
wire R18C28_GB10;
wire R1C47_S80;
wire VSS;
wire R6C17_GB10;
wire R1C1_N13;
wire R21C11_GB30;
wire R10C34_C5;
wire R12C12_GB10;
wire R13C5_GB60;
wire R26C43_GB10;
wire R22C24_GB30;
wire R5C30_GT10;
wire R18C43_GB50;
wire R1C28_C3;
wire R10C19_Q3;
wire R21C3_GBO0;
wire R12C32_GB50;
wire R28C43_B0;
wire R5C42_GBO0;
wire R14C32_GBO1;
wire R9C35_GB20;
wire R5C35_GB60;
wire R10C13_SEL0;
wire R28C28_D7;
wire R1C28_A3;
wire R18C45_GB70;
wire R23C6_GB40;
wire R28C22_S21;
wire R28C25_C4;
wire R17C40_GB00;
wire R20C5_SPINE19;
wire R5C12_GB30;
wire R18C9_GBO0;
wire R20C38_GB60;
wire R9C10_GT00;
wire R25C46_GBO1;
wire R1C28_Q4;
wire R10C34_N12;
wire R10C37_N11;
wire R25C7_GB00;
wire R4C37_GB20;
wire R23C22_GBO1;
wire R28C10_SEL0;
wire R14C13_GB40;
wire R2C36_GT00;
wire R21C2_GB70;
wire R6C29_GB40;
wire R20C37_GB70;
wire R10C10_X04;
wire R3C23_GB20;
wire R11C41_GB70;
wire R10C16_SEL2;
wire R10C16_S80;
wire R15C23_GB70;
wire R6C34_GB00;
wire R22C19_GB30;
wire R3C10_GT00;
wire R28C19_F4;
wire R26C19_GB30;
wire R15C5_GB70;
wire R28C34_S82;
wire R4C39_GBO0;
wire R4C20_GT00;
wire R2C24_GB40;
wire R16C11_GBO0;
wire R22C30_GB50;
wire R28C34_C7;
wire R16C24_GB20;
wire R10C13_F7;
wire R10C28_UNK127;
wire R28C19_C5;
wire R13C37_GB70;
wire R10C29_E13;
wire R8C24_GB70;
wire R20C14_GB20;
wire R29C28_X04;
wire R14C29_GBO1;
wire R28C43_D6;
wire R12C5_GB30;
wire R25C39_GB30;
wire R28C16_SEL4;
wire R28C22_Q1;
wire R26C2_GT10;
wire R28C19_Q4;
wire R28C16_SEL3;
wire R21C27_GB70;
wire R7C6_GB20;
wire R10C27_C1;
wire R28C46_A1;
wire R10C13_W12;
wire R10C34_D3;
wire R24C10_GB50;
wire R18C2_GB60;
wire R28C28_S81;
wire R13C23_GB20;
wire R17C46_GB60;
wire R7C25_GB70;
wire R21C13_GB50;
wire R6C10_GB70;
wire R18C11_GBO0;
wire R12C45_GB20;
wire R28C16_Q7;
wire R5C36_GB00;
wire R10C28_A0;
wire R22C13_GB40;
wire R22C8_GB60;
wire R28C22_N26;
wire R10C34_F6;
wire R28C43_W22;
wire R6C9_GB40;
wire R26C44_GBO1;
wire R16C35_GT00;
wire R5C39_GB20;
wire R1C32_D2;
wire R10C37_S23;
wire R23C4_GT10;
wire R11C16_GBO0;
wire R5C4_GB50;
wire R6C15_GB20;
wire R15C31_GT10;
wire R3C31_GB70;
wire R10C34_X08;
wire R17C23_GB40;
wire R10C31_C1;
wire R6C8_GT10;
wire R13C19_GB30;
wire R6C23_GB00;
wire R28C40_D5;
wire R18C4_GB40;
wire R14C33_GT10;
wire R10C7_CE2;
wire R14C11_GB00;
wire R12C16_GBO1;
wire R25C44_GB10;
wire R16C32_GB20;
wire R28C13_N26;
wire R28C25_X02;
wire R7C19_GB10;
wire R16C32_GBO1;
wire R15C15_GB40;
wire R1C28_A4;
wire R2C43_GBO0;
wire R13C14_GB10;
wire R24C17_GB50;
wire R8C45_GT00;
wire R29C28_D1;
wire R10C7_C3;
wire R15C17_GB50;
wire R2C6_GBO0;
wire R21C45_GT00;
wire R27C19_GB50;
wire R3C36_GT10;
wire R28C7_CLK0;
wire R28C10_N21;
wire R28C13_B2;
wire R26C12_GB50;
wire R17C20_GB70;
wire R3C41_GB50;
wire R25C15_GB60;
wire R28C43_S25;
wire R27C44_GB00;
wire R5C29_GT10;
wire R26C16_GBO0;
wire R16C37_GB00;
wire R1C1_A7;
wire R20C6_GB30;
wire R1C47_D5;
wire R16C18_GBO0;
wire R28C7_Q2;
wire R28C22_D6;
wire R10C16_D4;
wire R10C25_X05;
wire R6C42_GB60;
wire R4C10_GB30;
wire R8C21_GBO0;
wire R15C39_GB50;
wire R8C18_GB50;
wire R2C34_GB20;
wire R6C3_GB00;
wire R28C4_B6;
wire R28C37_CLK0;
wire R3C15_GB10;
wire R10C29_UNK121;
wire R28C31_SEL2;
wire R7C8_GB10;
wire R11C4_GBO1;
wire R14C33_GT00;
wire R22C26_GB10;
wire R11C42_GB20;
wire R10C10_X07;
wire R10C31_N10;
wire R3C36_GB20;
wire R14C31_GB50;
wire R28C10_W13;
wire R13C2_GB30;
wire R17C9_GB00;
wire R24C30_GB20;
wire R22C22_GT10;
wire R22C33_GT00;
wire R24C9_GB10;
wire R14C7_GB70;
wire R26C42_GBO1;
wire R20C14_GBO1;
wire R12C38_GB70;
wire R7C35_GT10;
wire R16C17_GB50;
wire R7C21_GB00;
wire R10C25_S21;
wire R22C39_GB60;
wire R11C13_GBO1;
wire R15C19_GB60;
wire R18C18_GB00;
wire R7C14_GT00;
wire R5C29_GB50;
wire R23C45_GB60;
wire R17C10_GB40;
wire R26C19_GB70;
wire R5C3_GBO0;
wire R3C3_GB20;
wire R27C7_GBO1;
wire R13C36_GB20;
wire R1C32_C7;
wire R10C25_LSR1;
wire R28C28_X02;
wire R28C37_N22;
wire R28C46_SEL0;
wire R25C7_GB50;
wire R10C28_A4;
wire R3C28_GB00;
wire R1C28_S23;
wire R5C17_GBO0;
wire R17C14_GB60;
wire R20C34_GB60;
wire R10C28_D3;
wire R11C7_GB70;
wire R6C5_GB20;
wire R16C23_GT00;
wire R2C31_GT10;
wire R8C34_GBO0;
wire R12C34_GB30;
wire R21C9_GB40;
wire R11C4_GBO0;
wire R5C34_GBO1;
wire R22C28_GT00;
wire R5C36_GT00;
wire R20C41_GB50;
wire R9C20_GB60;
wire R3C20_GB20;
wire R5C30_GB30;
wire R28C25_S80;
wire R26C16_GB30;
wire R28C7_E10;
wire R7C6_GB70;
wire R20C17_GT10;
wire R9C35_GB60;
wire R26C4_GB30;
wire R14C2_GT00;
wire R12C14_GB40;
wire R23C2_GB30;
wire R27C19_GB70;
wire R14C11_GB30;
wire R6C31_GB70;
wire R10C43_S13;
wire R22C42_GB70;
wire R28C4_Q2;
wire R8C4_GBO0;
wire R29C28_X02;
wire R10C30_F7;
wire R4C28_GB40;
wire R24C3_GT10;
wire R10C37_E22;
wire R21C24_GBO1;
wire R10C16_X04;
wire R21C45_GB30;
wire R28C22_W82;
wire R23C22_GT10;
wire R11C35_GBO0;
wire R4C33_GT00;
wire R9C21_GB60;
wire R1C28_N24;
wire R4C15_GB70;
wire R10C25_B5;
wire R17C41_GB20;
wire R10C16_F7;
wire R28C34_A0;
wire R26C8_GT00;
wire R20C6_GB10;
wire R2C34_GB00;
wire R22C37_GBO0;
wire R10C25_SEL5;
wire R17C8_GB20;
wire R7C33_GB40;
wire R25C35_GT00;
wire R10C30_X01;
wire R10C31_S12;
wire R8C38_GB00;
wire R20C20_SPINE20;
wire R10C34_CLK0;
wire R28C25_S12;
wire R22C8_GT00;
wire R28C13_B6;
wire R26C8_GB40;
wire R23C16_GT00;
wire R27C7_GB20;
wire R23C20_GB20;
wire R24C3_GB30;
wire R9C36_GB20;
wire R28C19_N20;
wire R13C4_GB00;
wire R27C6_GT00;
wire R13C45_GB70;
wire R28C46_E23;
wire R2C4_GB50;
wire R28C46_E22;
wire R11C30_GB40;
wire R8C44_GBO1;
wire R1C28_D1;
wire R27C22_GB20;
wire R17C30_GBO0;
wire R27C16_GB50;
wire R8C22_GBO0;
wire R22C46_GB70;
wire R7C5_GBO1;
wire R24C34_GB40;
wire R28C10_C4;
wire R20C20_GBO0;
wire R12C11_GT00;
wire R25C17_GB30;
wire R26C10_GB60;
wire R10C10_D5;
wire R14C9_GBO0;
wire R5C43_GBO0;
wire R16C4_GB70;
wire R10C26_D5;
wire R10C25_S80;
wire R7C18_GBO0;
wire R8C22_GT10;
wire R28C22_S13;
wire R28C10_C1;
wire R12C3_GT00;
wire R18C2_GB70;
wire R13C24_GBO1;
wire R22C31_GB50;
wire R6C44_GB20;
wire R27C22_GB70;
wire R24C31_GB20;
wire R16C5_GB10;
wire R28C34_S11;
wire R22C44_GB40;
wire R14C8_GT00;
wire R3C16_GB40;
wire R20C26_GB60;
wire R11C4_GB50;
wire R22C42_GB60;
wire R18C24_GB40;
wire R3C15_GT10;
wire R16C40_GB40;
wire R12C35_GBO1;
wire R10C40_D6;
wire R25C9_GB30;
wire R13C4_GT00;
wire R14C36_GB60;
wire R16C29_GT10;
wire R22C32_GBO0;
wire R10C37_S12;
wire R10C29_W25;
wire R4C19_GB40;
wire R8C4_GB00;
wire R4C29_GB30;
wire R16C14_GT00;
wire R8C35_GB60;
wire R15C13_GBO1;
wire R28C7_EW20;
wire R3C41_GB70;
wire R7C9_GB60;
wire R8C22_GB00;
wire R26C30_GBO0;
wire R10C19_D6;
wire R10C31_S26;
wire R10C22_F2;
wire R28C40_B2;
wire R7C38_GT00;
wire R23C6_GBO0;
wire R21C42_GB50;
wire R28C40_D1;
wire R25C5_GB60;
wire R26C11_GB10;
wire R10C27_A5;
wire R28C37_Q5;
wire R12C5_GB50;
wire R1C47_W13;
wire R3C35_GB20;
wire R17C45_GB20;
wire R20C16_GB70;
wire R28C22_CLK0;
wire R10C28_E80;
wire R8C45_GBO0;
wire R3C18_GB00;
wire R24C21_GBO0;
wire R14C41_GB20;
wire R27C34_GB60;
wire R1C47_W23;
wire R10C10_F1;
wire R10C19_SEL0;
wire R11C20_GB50;
wire R23C12_GB10;
wire R9C7_GT10;
wire R10C34_EW20;
wire R26C39_GB20;
wire R6C22_GB60;
wire R10C37_W11;
wire R28C46_S82;
wire R21C38_GB20;
wire R28C28_S83;
wire R27C11_GT10;
wire R28C34_N24;
wire R27C46_GB10;
wire R23C8_GB60;
wire R17C27_GB10;
wire R4C6_GB30;
wire R25C33_GB20;
wire R26C39_GT00;
wire R16C14_GB60;
wire R28C7_E83;
wire R12C13_GB60;
wire R11C39_GT10;
wire R21C32_GB00;
wire R27C7_GB00;
wire R25C26_GBO0;
wire R23C9_GB40;
wire R4C7_GB30;
wire R10C43_D6;
wire R24C28_GT00;
wire R13C38_GT00;
wire R5C20_GBO1;
wire R8C31_GB10;
wire R10C7_S13;
wire R28C46_LSR2;
wire R10C25_SEL0;
wire R10C22_E25;
wire R26C13_GBO0;
wire R10C31_N26;
wire R28C4_F7;
wire R24C23_GT10;
wire R3C27_GBO1;
wire R16C19_GB20;
wire R26C5_GB10;
wire R16C23_GB10;
wire R10C34_E80;
wire R10C43_S23;
wire R2C4_GB40;
wire R13C5_GB40;
wire R5C22_GB10;
wire R12C20_GBO1;
wire R20C44_GB10;
wire R9C39_GB20;
wire R3C31_GT10;
wire R10C29_UNK126;
wire R13C10_GB40;
wire R25C7_GB60;
wire R23C32_GB60;
wire R14C3_GBO0;
wire R10C16_SEL0;
wire R28C31_EW20;
wire R18C27_GB20;
wire R28C25_X07;
wire R23C9_GB00;
wire R25C39_GB10;
wire R17C29_GB20;
wire R15C35_GB30;
wire R14C27_GT10;
wire R18C6_GBO0;
wire R1C28_F4;
wire R10C34_SEL4;
wire R10C40_W20;
wire R10C37_S21;
wire R25C15_GB30;
wire R21C40_GB50;
wire R23C3_GB20;
wire R11C16_GB30;
wire R25C8_GB60;
wire R10C34_W11;
wire R16C21_GB60;
wire R8C45_GB20;
wire R12C9_GB50;
wire R8C29_GB10;
wire R1C32_C2;
wire R15C38_GT00;
wire R1C1_A6;
wire R10C29_N27;
wire R7C33_GBO0;
wire R1C1_B4;
wire R10C16_D5;
wire R13C19_GB40;
wire R11C9_GB50;
wire R1C32_S10;
wire R10C13_Q2;
wire R10C25_S12;
wire R28C31_W10;
wire R12C21_GB30;
wire R9C17_GB60;
wire R6C43_GB30;
wire R9C23_GB00;
wire R7C15_GB50;
wire R17C17_GBO1;
wire R6C6_GB60;
wire R28C7_F7;
wire R18C14_GT10;
wire R20C21_GB00;
wire R15C45_GB70;
wire R10C10_SEL5;
wire R28C25_W83;
wire R14C38_GB40;
wire R22C11_GT00;
wire R18C13_GB50;
wire R24C43_GBO0;
wire R10C7_D7;
wire R7C17_GBO1;
wire R26C22_GT00;
wire R28C28_Q5;
wire R15C14_GB50;
wire R10C43_A4;
wire R28C22_N25;
wire R23C44_GB50;
wire R10C30_LSR2;
wire R2C12_GB70;
wire R23C13_GBO1;
wire R10C16_E26;
wire R14C30_GT10;
wire R3C14_GB10;
wire R9C9_GB70;
wire R25C25_GB40;
wire R2C38_GB00;
wire R1C47_N13;
wire R10C29_W26;
wire R15C23_GB60;
wire R24C17_GB10;
wire R21C27_GB60;
wire R3C12_GB60;
wire R22C44_GB50;
wire R10C31_B5;
wire R28C7_F5;
wire R21C34_GB00;
wire R28C10_Q1;
wire R3C32_GB10;
wire R22C34_GB10;
wire R12C11_GB00;
wire R3C37_GB30;
wire R8C15_GB00;
wire R9C40_GT10;
wire R16C13_GB60;
wire R27C20_GB20;
wire R10C29_B5;
wire R16C7_GB10;
wire R3C35_GB30;
wire R7C20_GT00;
wire R5C38_GB10;
wire R8C8_GB40;
wire R3C22_GB50;
wire R10C34_SEL0;
wire R28C4_C4;
wire R12C12_GT10;
wire R5C4_GB30;
wire R18C8_GB00;
wire R24C16_GB30;
wire R1C32_EW10;
wire R2C34_SPINE2;
wire R3C23_GT00;
wire R24C27_GB10;
wire R28C10_Q0;
wire R28C22_D5;
wire R10C31_X08;
wire R28C10_C0;
wire R23C25_GT10;
wire R7C11_GB50;
wire R10C26_S11;
wire R8C27_GB40;
wire R4C42_GB40;
wire R1C47_LSR1;
wire R13C8_GB20;
wire R21C35_GB70;
wire R28C7_A4;
wire R12C4_GB70;
wire R10C28_N26;
wire R25C30_GB00;
wire R10C28_SPINE20;
wire R28C4_SEL7;
wire R20C36_GB60;
wire R4C24_GB40;
wire R11C38_GB00;
wire R22C36_GBO1;
wire R10C25_N82;
wire R10C26_E20;
wire R10C27_N24;
wire R27C18_GB00;
wire R21C14_GT10;
wire R8C21_GB50;
wire R22C25_GB10;
wire R26C37_GT10;
wire R22C13_GBO0;
wire R16C23_GB30;
wire R20C1_GBO1;
wire R10C37_C4;
wire R6C9_GT10;
wire R10C37_SN20;
wire R8C35_GB20;
wire R13C31_GBO0;
wire R13C37_GT00;
wire R5C9_GB30;
wire R28C40_S13;
wire R17C28_GB60;
wire R12C37_GB20;
wire R23C33_GBO0;
wire R15C38_GB60;
wire R16C36_GB60;
wire R28C40_LSR2;
wire R14C39_GB30;
wire R10C25_F7;
wire R10C31_N80;
wire R16C10_GB70;
wire R5C44_GB60;
wire R20C16_GT10;
wire R15C5_GT10;
wire R26C17_GB00;
wire R4C6_GB40;
wire R20C23_GT10;
wire R14C44_GT00;
wire R15C21_GB20;
wire R12C21_GB50;
wire R13C1_GT10;
wire R26C29_GB50;
wire R2C39_GBO1;
wire R14C42_GB00;
wire R9C22_GB20;
wire R4C1_GBO1;
wire R5C24_GB70;
wire R11C19_GB30;
wire R27C43_GB70;
wire R10C19_SEL7;
wire R10C13_Q3;
wire R2C16_GB00;
wire R25C17_GBO0;
wire R10C28_E27;
wire R23C29_GBO1;
wire R18C40_GB00;
wire R10C40_SN10;
wire R28C34_S12;
wire R28C43_E23;
wire R12C15_GB00;
wire R5C40_GB70;
wire R11C1_GBO1;
wire R5C29_GB00;
wire R28C34_CLK0;
wire R25C20_GT10;
wire R13C35_GBO1;
wire R3C19_GB30;
wire R14C21_GBO0;
wire R3C33_GB00;
wire R6C34_GB10;
wire R26C35_GB50;
wire R28C22_X07;
wire R22C15_GBO0;
wire R14C34_GT10;
wire R4C38_GBO0;
wire R5C13_GB10;
wire R9C15_GB20;
wire R28C19_C3;
wire R10C25_W13;
wire R6C44_GB60;
wire R10C19_W24;
wire R5C19_GB10;
wire R5C4_GB70;
wire R18C37_GB20;
wire R11C28_GB10;
wire R28C13_S20;
wire R27C11_GB20;
wire R8C27_GB20;
wire R26C32_GB40;
wire R8C25_GB50;
wire R10C28_UNK123;
wire R11C38_GT10;
wire R28C4_N22;
wire R28C31_N11;
wire R18C30_GT00;
wire R2C18_GB70;
wire R14C16_GBO0;
wire R2C41_GBO1;
wire R8C25_GB70;
wire R22C30_GB70;
wire R28C25_SEL6;
wire R28C46_D6;
wire R17C34_GB70;
wire R8C2_GBO1;
wire R13C25_GB50;
wire R7C29_GB10;
wire R22C24_GT00;
wire R5C11_GB60;
wire R20C42_GB10;
wire R24C21_GT10;
wire R28C37_S26;
wire R21C23_GT00;
wire R27C28_GB20;
wire R10C29_E24;
wire R12C34_GB40;
wire R10C27_E10;
wire R11C18_GB30;
wire R27C18_GT10;
wire R25C18_GB30;
wire R3C5_GT10;
wire R21C22_GB30;
wire R25C28_GB40;
wire R16C42_GB10;
wire R11C34_GB50;
wire R1C32_SEL0;
wire R10C19_Q0;
wire R10C19_F5;
wire R28C7_S82;
wire R1C47_CE0;
wire R10C30_E82;
wire R24C12_GB50;
wire R4C3_GB40;
wire R16C20_GB10;
wire R24C39_GB50;
wire R18C19_GB20;
wire R12C9_GB00;
wire R10C10_W11;
wire R9C46_GB70;
wire R1C47_F0;
wire R11C37_GB00;
wire R15C5_GB40;
wire R18C41_GB20;
wire R4C7_GBO0;
wire R10C16_F4;
wire R10C28_B5;
wire R18C44_GB40;
wire R21C10_GB20;
wire R26C44_GB70;
wire R10C31_CE2;
wire R28C34_SEL0;
wire R11C25_GB00;
wire R5C44_GB20;
wire R8C46_GT00;
wire R2C24_GT00;
wire R3C21_GB20;
wire R24C8_GB10;
wire R28C22_SN20;
wire R27C45_GT10;
wire R21C6_GB40;
wire R11C12_GB60;
wire R18C43_GB00;
wire R1C47_S26;
wire R1C32_X01;
wire R10C27_W26;
wire R22C24_GBO1;
wire R6C46_GB50;
wire R27C12_GB70;
wire R7C4_GB70;
wire R27C15_GB40;
wire R5C36_GB40;
wire R1C1_B7;
wire R28C13_SN20;
wire R28C4_C2;
wire R2C19_GB10;
wire R7C28_GB70;
wire R22C9_GB30;
wire R21C6_GT00;
wire R7C22_GB40;
wire R27C19_GB20;
wire R10C40_F7;
wire R6C29_GB10;
wire R23C19_GB70;
wire R16C30_GT10;
wire R12C15_GB50;
wire R8C32_GB20;
wire R28C10_X05;
wire R3C2_GB50;
wire R23C37_GB20;
wire R10C43_N24;
wire R8C9_GB50;
wire R4C43_GB10;
wire R3C2_GB20;
wire R8C38_GB40;
wire R1C32_SN20;
wire R10C25_E21;
wire R14C27_GB30;
wire R10C43_C1;
wire R7C31_GB40;
wire R13C34_GB20;
wire R21C6_GB10;
wire R13C20_GB40;
wire R29C28_SEL6;
wire R9C7_GT00;
wire R5C42_GB40;
wire R28C25_E12;
wire R1C47_N83;
wire R24C7_GBO0;
wire R20C29_GT10;
wire R11C38_GB30;
wire R24C36_GT00;
wire R10C34_S82;
wire R5C20_GT10;
wire R25C43_GBO1;
wire R28C16_C4;
wire R13C27_GT10;
wire R29C28_N23;
wire R5C25_GBO0;
wire R28C43_E80;
wire R12C11_GB50;
wire R10C31_LSR0;
wire R7C35_GBO0;
wire R23C5_GT10;
wire R9C11_GB60;
wire R23C6_GB50;
wire R27C35_GB10;
wire R5C23_GB40;
wire R25C17_GB20;
wire R21C43_GB10;
wire R11C44_GT00;
wire R4C40_GT00;
wire R10C27_D3;
wire R20C40_GBO1;
wire R24C12_GT10;
wire R24C27_GT00;
wire R4C7_GB70;
wire R4C14_GB40;
wire R24C17_GB20;
wire R7C18_GT10;
wire R27C16_GB70;
wire R11C1_GT10;
wire R12C9_GT10;
wire R3C8_GB10;
wire R9C36_GB70;
wire R1C28_E80;
wire R18C11_GB10;
wire R10C26_Q5;
wire R10C28_SEL6;
wire R8C34_GT00;
wire R28C37_S11;
wire R25C41_GB40;
wire R6C25_GB40;
wire R7C35_GB30;
wire R20C38_GT00;
wire R4C37_GBO1;
wire R6C40_GB10;
wire R2C26_GB20;
wire R25C37_GBO1;
wire R4C9_GT10;
wire R11C19_GB60;
wire R12C14_GT10;
wire R10C34_E25;
wire R13C41_GB10;
wire R24C15_GB70;
wire R24C4_GB40;
wire R8C23_GB10;
wire R13C40_GT10;
wire R24C9_GB00;
wire R12C7_GBO0;
wire R22C16_GBO1;
wire R21C10_GB50;
wire R1C47_E27;
wire R10C30_Q7;
wire R29C28_B4;
wire R26C22_GBO1;
wire R28C43_SN10;
wire R21C36_GB20;
wire R24C35_GBO0;
wire R4C4_GB30;
wire R14C43_GBO0;
wire R25C44_GB70;
wire R7C10_GB20;
wire R23C20_GT00;
wire R14C15_GBO1;
wire R28C10_D6;
wire R27C45_GB20;
wire R27C38_GB40;
wire R10C30_Q2;
wire R4C2_GBO1;
wire R8C7_GB40;
wire R10C26_EW20;
wire R2C33_GB00;
wire R10C28_SPINE19;
wire R28C28_SEL7;
wire R10C25_E23;
wire R27C42_GB60;
wire R25C21_GB60;
wire R25C46_GT00;
wire R5C16_GBO1;
wire R13C7_GT00;
wire R14C25_GB10;
wire R2C3_GT00;
wire R26C46_GT10;
wire R14C15_GB70;
wire R13C13_GBO1;
wire R4C20_GB50;
wire R6C19_GB30;
wire R25C31_GB30;
wire R28C10_B3;
wire R20C11_GB30;
wire R29C28_S83;
wire R27C19_GBO0;
wire R15C37_GBO1;
wire R28C25_E20;
wire R20C3_GB50;
wire R20C25_GB60;
wire R2C20_GBO0;
wire R12C29_GB40;
wire R6C10_GT00;
wire R4C17_GBO1;
wire R22C16_GB10;
wire R20C21_GT00;
wire R9C35_GT00;
wire R6C25_GB00;
wire R3C16_GB30;
wire R10C13_D7;
wire R22C2_GT00;
wire R10C19_B5;
wire R28C28_E12;
wire R10C25_Q6;
wire R1C28_SEL6;
wire R4C45_GB00;
wire R25C40_GBO0;
wire R11C34_GB10;
wire R10C10_W10;
wire R21C7_GB60;
wire R29C28_W11;
wire R20C14_GB10;
wire R16C8_GBO0;
wire R11C11_GB20;
wire R10C31_SEL0;
wire R3C37_GT00;
wire R27C30_GB60;
wire R22C33_GBO0;
wire R2C44_GBO0;
wire R21C2_GB50;
wire R10C40_N81;
wire R10C7_Q4;
wire R25C2_GB30;
wire R26C24_GB20;
wire R10C16_B6;
wire R7C45_GB20;
wire R21C30_GT00;
wire R9C5_GB30;
wire R21C29_GB50;
wire R20C24_GB20;
wire R12C23_GBO1;
wire R10C28_E22;
wire R6C32_GB50;
wire R10C10_E11;
wire R1C28_F7;
wire R28C4_W11;
wire R10C16_CLK1;
wire R10C40_B5;
wire R2C41_GB20;
wire R4C22_GB60;
wire R12C19_GB50;
wire R9C41_GB10;
wire R11C11_GB40;
wire R12C6_GB50;
wire R10C13_LSR2;
wire R18C12_GBO1;
wire R10C16_S82;
wire R28C34_N21;
wire R28C40_SEL7;
wire R12C29_GB10;
wire R10C30_F5;
wire R10C40_B3;
wire R28C34_E83;
wire R18C11_GT10;
wire R3C8_GB70;
wire R15C32_GBO0;
wire R10C10_W13;
wire R7C43_GB70;
wire R28C40_W20;
wire R14C13_GB30;
wire R29C28_S80;
wire R12C38_GB00;
wire R16C34_GB00;
wire R12C21_GBO0;
wire R18C25_GB40;
wire R25C16_GT00;
wire R3C20_GB70;
wire R20C5_GB30;
wire R18C38_GBO0;
wire R28C4_B4;
wire R17C23_GB30;
wire R3C10_GT10;
wire R5C23_GBO1;
wire R26C21_GB70;
wire R20C33_GB40;
wire R3C10_GB30;
wire R11C27_GB20;
wire R27C46_GB30;
wire R17C32_GT10;
wire R10C25_S25;
wire R7C24_GB70;
wire R10C27_LSR0;
wire R2C12_GBO1;
wire R13C31_GT00;
wire R27C19_GT10;
wire R6C11_GB20;
wire R10C19_LSR0;
wire R9C43_GB30;
wire R16C32_GT00;
wire R7C27_GB60;
wire R10C43_A2;
wire R2C9_GT00;
wire R3C35_GT10;
wire R8C15_GB40;
wire R3C15_GBO1;
wire R16C13_GT10;
wire R28C37_E13;
wire R17C5_GB30;
wire R20C20_GT10;
wire R25C39_GB60;
wire R7C40_GB00;
wire R18C11_GBO1;
wire R7C44_GB30;
wire R15C32_GB70;
wire R5C21_GBO1;
wire R16C5_GB40;
wire R6C25_GB10;
wire R22C9_GB20;
wire R18C35_GB40;
wire R10C30_EW10;
wire R28C7_S23;
wire R28C40_A0;
wire R9C42_GBO1;
wire R27C42_GB00;
wire R12C22_GB40;
wire R13C3_GB40;
wire R9C44_GBO0;
wire R28C43_A3;
wire R10C43_S26;
wire R17C14_GB30;
wire R4C28_GB50;
wire R26C39_GBO1;
wire R1C47_CE1;
wire R17C39_GB70;
wire R10C7_F3;
wire R28C25_B6;
wire R18C10_GB60;
wire R28C46_E12;
wire R5C9_GBO1;
wire R22C19_GB70;
wire R7C33_GB10;
wire R10C27_A3;
wire R10C28_N80;
wire R10C29_W24;
wire R28C4_S26;
wire R27C3_GB60;
wire R3C24_GB50;
wire R10C10_Q2;
wire R11C21_GB30;
wire R10C7_D4;
wire R10C40_Q7;
wire R9C43_GB00;
wire R1C1_A1;
wire R10C28_F6;
wire R29C28_Q1;
wire R7C40_GB40;
wire R10C25_W23;
wire R27C16_GT10;
wire R4C21_GBO0;
wire R22C34_GB30;
wire R10C13_S26;
wire R12C10_GB20;
wire R6C27_GB20;
wire R28C25_Q6;
wire R16C7_GB60;
wire R28C40_Q1;
wire R3C41_GB30;
wire R28C7_N22;
wire R28C43_LSR0;
wire R27C28_GT10;
wire R2C12_GB50;
wire R22C17_GB20;
wire R8C10_GB00;
wire R2C22_GB20;
wire R10C43_W25;
wire R21C31_GT10;
wire R28C7_X05;
wire R15C18_GB10;
wire R17C18_GB30;
wire R27C3_GB70;
wire R21C46_GB00;
wire R16C37_GB20;
wire R7C7_GB30;
wire R8C29_GB00;
wire R1C1_N22;
wire R14C18_GB50;
wire R1C28_E81;
wire R10C34_C0;
wire R10C16_F2;
wire R11C45_GB20;
wire R13C4_GT10;
wire R16C35_GB20;
wire R28C40_CLK0;
wire R27C37_GB50;
wire R21C43_GB50;
wire R1C47_SEL0;
wire R28C31_C6;
wire R10C34_W83;
wire R1C32_W25;
wire R7C5_GB30;
wire R8C7_GBO0;
wire R5C40_GBO0;
wire R5C40_GB60;
wire R26C26_GT10;
wire R15C31_GB10;
wire R6C3_GBO0;
wire R4C22_GB50;
wire R15C31_GB50;
wire R10C10_X06;
wire R10C28_LSR2;
wire R28C34_B6;
wire R21C21_GB20;
wire R10C31_A6;
wire R6C2_GB40;
wire R28C19_CE1;
wire R11C22_GBO1;
wire R27C45_GB10;
wire R7C10_GBO1;
wire R21C7_GB20;
wire R10C7_N21;
wire R10C7_E25;
wire R21C46_GBO0;
wire R10C37_F0;
wire R28C25_X04;
wire R10C25_A1;
wire R18C12_GT00;
wire R3C36_GB00;
wire R4C25_GB00;
wire R22C36_GB70;
wire R7C41_GB00;
wire R6C5_GB60;
wire R13C6_GBO0;
wire R21C7_GB50;
wire R11C45_GBO0;
wire R24C26_GT00;
wire R20C8_GB50;
wire R10C31_CE0;
wire R28C13_CE0;
wire R18C22_GT00;
wire R27C46_GBO1;
wire R28C22_X01;
wire R8C7_GT10;
wire R22C17_GB60;
wire R15C25_GBO1;
wire R10C31_W13;
wire R24C38_GB30;
wire R6C22_GB10;
wire R20C12_GT10;
wire R9C17_GB20;
wire R18C26_GB50;
wire R2C18_GB30;
wire R14C27_GB20;
wire R24C6_GT10;
wire R5C13_GB20;
wire R2C3_GB70;
wire R7C5_GB70;
wire R6C29_GB70;
wire R16C39_GB30;
wire R23C16_GB60;
wire R28C7_C7;
wire R28C34_C0;
wire R14C43_GT10;
wire R28C34_F2;
wire R12C22_GBO1;
wire R17C7_GB40;
wire R2C42_GB60;
wire R4C22_GB10;
wire R7C45_GB50;
wire R26C17_GB10;
wire R9C16_GBO1;
wire R8C20_GB50;
wire R15C18_GT00;
wire R13C14_GB00;
wire R28C10_B2;
wire R18C30_GB20;
wire R29C28_LSR1;
wire R16C37_GB50;
wire R26C44_GB20;
wire R5C13_GB40;
wire R10C37_N10;
wire R11C43_GB50;
wire R8C24_GBO0;
wire R27C12_GB40;
wire R4C16_GB60;
wire R9C38_GB60;
wire R18C45_GB00;
wire R14C22_GB70;
wire R25C45_GB10;
wire R26C41_GT00;
wire R17C24_GBO0;
wire R6C30_GB60;
wire R13C38_GB70;
wire R2C19_GB70;
wire R13C30_GB30;
wire R5C44_GBO0;
wire R27C32_GB50;
wire R1C1_CE2;
wire R16C18_GB40;
wire R10C13_Q6;
wire R2C38_GB60;
wire R28C22_N80;
wire R10C29_N23;
wire R25C27_GB10;
wire R17C11_GBO0;
wire R15C22_GB10;
wire R24C45_GB20;
wire R14C32_GB40;
wire R10C29_N10;
wire R28C28_S21;
wire R8C44_GBO0;
wire R28C46_F7;
wire R25C2_GB00;
wire R15C39_GBO1;
wire R17C41_GBO1;
wire R16C4_GT00;
wire R28C25_A4;
wire R28C40_S24;
wire R16C16_GT10;
wire R27C42_GT10;
wire R2C39_GB30;
wire R22C35_GBO1;
wire R1C28_CE1;
wire R4C11_GB60;
wire R10C28_B1;
wire R14C26_GB70;
wire R4C22_GT10;
wire R13C39_GB70;
wire R10C34_B0;
wire R28C7_W10;
wire R22C16_GB60;
wire R6C39_GBO1;
wire R22C5_GB70;
wire R3C26_GB00;
wire R11C2_GB40;
wire R4C13_GBO1;
wire R24C30_GB70;
wire R22C38_GB70;
wire R24C10_GBO1;
wire R3C27_GBO0;
wire R10C40_E81;
wire R7C28_GB40;
wire R2C6_GB60;
wire R27C16_GBO0;
wire R24C24_GBO0;
wire R7C46_GBO1;
wire R10C26_W12;
wire R10C30_W21;
wire R5C18_GBO0;
wire R10C34_N21;
wire R28C13_CE2;
wire R13C25_GB20;
wire R22C29_GB70;
wire R4C2_GT00;
wire R15C14_GB70;
wire R3C11_GB30;
wire R28C46_W12;
wire R25C26_GB60;
wire R8C10_GB60;
wire R27C24_GB20;
wire R23C44_GT00;
wire R12C38_GB60;
wire R9C38_GB30;
wire R28C13_N23;
wire R26C23_GT00;
wire R17C16_GBO1;
wire R27C8_GB00;
wire R23C22_GB50;
wire R28C40_N80;
wire R10C43_A3;
wire R1C28_S12;
wire R7C3_GB40;
wire R28C46_SEL1;
wire R5C45_GT00;
wire R25C4_GB40;
wire R21C16_GB40;
wire R9C36_GB10;
wire R28C4_D4;
wire R18C24_GB00;
wire R8C37_GB20;
wire R4C22_GB00;
wire R22C45_GB70;
wire R22C32_GBO1;
wire R25C27_GT00;
wire R28C28_D5;
wire R27C41_GB40;
wire R12C43_GB60;
wire R10C7_E24;
wire R20C7_GB00;
wire R27C10_GT10;
wire R3C21_GT10;
wire R25C38_GB20;
wire R13C44_GB50;
wire R28C16_E13;
wire R4C2_GB20;
wire R2C33_GT10;
wire R26C3_GB40;
wire R18C4_GB60;
wire R28C28_A6;
wire R24C15_GT00;
wire R3C15_GT00;
wire R15C10_GB40;
wire R22C12_GB40;
wire R28C7_N23;
wire R28C19_E12;
wire R20C6_SPINE18;
wire R27C38_GB30;
wire R28C37_SEL2;
wire R11C34_GBO0;
wire R6C39_GB00;
wire R4C8_GB00;
wire R25C45_GB30;
wire R28C16_D2;
wire R22C37_GBO1;
wire R14C17_GBO1;
wire R10C16_CE0;
wire R24C44_GT00;
wire R6C6_GB00;
wire R16C21_GB10;
wire R23C21_GB20;
wire R27C25_GB70;
wire R28C16_A5;
wire R10C29_S22;
wire R6C26_GB50;
wire R11C24_GB10;
wire R24C27_GB00;
wire R28C25_E23;
wire R26C24_GB00;
wire R9C20_GB30;
wire R25C15_GBO1;
wire R27C26_GT10;
wire R23C45_GB20;
wire R1C32_LSR0;
wire R9C24_GB40;
wire R1C1_S24;
wire R28C7_SN10;
wire R23C27_GB50;
wire R15C35_GB00;
wire R9C38_GB70;
wire R10C27_N82;
wire R10C30_N81;
wire R28C10_EW10;
wire R20C17_GBO0;
wire R26C38_GB00;
wire R12C40_GBO0;
wire R21C31_GB10;
wire R18C36_GBO0;
wire R10C34_S20;
wire R21C12_GT10;
wire R28C16_F1;
wire R16C2_GBO0;
wire R20C7_GBO0;
wire R22C29_GT00;
wire R25C12_GBO1;
wire R28C46_N81;
wire R16C27_GB00;
wire R3C42_GBO0;
wire R6C30_GT00;
wire R11C21_GBO1;
wire R3C41_GB00;
wire R29C28_C5;
wire R18C42_GB30;
wire R20C40_GT10;
wire R16C18_GB60;
wire R10C26_S21;
wire R10C27_Q3;
wire R28C31_N82;
wire R17C24_GB60;
wire R24C36_GBO1;
wire R10C7_E21;
wire R6C20_GT00;
wire R4C44_GB10;
wire R23C5_GB00;
wire R6C22_GT10;
wire R13C32_GB50;
wire R10C27_B3;
wire R7C39_GB50;
wire R16C19_GBO1;
wire R22C38_GBO0;
wire R15C20_GB10;
wire R8C39_GB50;
wire R6C16_GB20;
wire R5C7_GB10;
wire R13C37_GB00;
wire R10C7_B3;
wire R26C37_GB50;
wire R28C40_CE2;
wire R20C40_GB10;
wire R28C16_W23;
wire R2C25_GB10;
wire R4C19_GB50;
wire R15C16_GB10;
wire R28C40_LSR0;
wire R16C26_GT00;
wire R22C20_GT10;
wire R5C27_GB40;
wire R1C32_SEL2;
wire R23C14_GB20;
wire R23C31_GB30;
wire R15C26_GB10;
wire R10C28_W23;
wire R25C23_GB60;
wire R18C5_GBO1;
wire R20C22_GT10;
wire R21C38_GB60;
wire R28C13_EW20;
wire R26C45_GB60;
wire R14C44_GB60;
wire R10C34_A7;
wire R28C43_Q0;
wire R2C22_GB10;
wire R22C11_GBO1;
wire R10C43_SEL2;
wire R20C11_SPINE21;
wire R8C2_GBO0;
wire R28C31_SEL0;
wire R3C14_GT10;
wire R11C19_GBO1;
wire R5C15_GB10;
wire R5C46_GB30;
wire R4C45_GB60;
wire R12C32_GB30;
wire R23C5_GBO0;
wire R13C33_GB50;
wire R1C47_W81;
wire R10C28_S11;
wire R5C29_GB20;
wire R5C42_GB00;
wire R22C18_GBO1;
wire R26C30_GB70;
wire R5C9_GB20;
wire R13C41_GB20;
wire R28C31_E22;
wire R1C28_C6;
wire R10C16_A6;
wire R13C33_GB20;
wire R22C9_GBO0;
wire R1C47_B4;
wire R28C37_S27;
wire R9C8_GT00;
wire R10C25_SEL7;
wire R12C34_GBO1;
wire R21C42_GB30;
wire R22C45_GB00;
wire R26C15_GB10;
wire R14C14_GB10;
wire R10C34_SEL3;
wire R4C4_GB40;
wire R10C13_S10;
wire R4C37_GB10;
wire R18C25_GT10;
wire R7C38_GB10;
wire R24C29_GB10;
wire R17C15_GB50;
wire R26C39_GB10;
wire R27C32_GB40;
wire R1C47_S21;
wire R5C11_GB10;
wire R23C31_GB50;
wire R27C44_GT00;
wire R23C33_GT10;
wire R10C22_N23;
wire R15C29_GB70;
wire R4C31_GB60;
wire R10C34_E24;
wire R17C39_GB50;
wire R10C31_B7;
wire R6C15_GB10;
wire R21C3_GBO1;
wire R5C39_GB60;
wire R23C32_GB40;
wire R7C11_GB60;
wire R10C19_N82;
wire R10C37_Q2;
wire R28C46_W24;
wire R10C19_W20;
wire R26C30_GB20;
wire R28C37_W25;
wire R4C23_GBO1;
wire R28C19_A1;
wire R3C18_GB70;
wire R26C36_GB40;
wire R9C28_GB50;
wire R27C36_GT10;
wire R9C11_GB00;
wire R10C40_Q4;
wire R5C36_GB10;
wire R10C10_D6;
wire R28C4_F6;
wire R8C24_GB00;
wire R20C38_GB10;
wire R11C17_GB60;
wire R27C17_GB20;
wire R3C37_GB50;
wire R28C31_S83;
wire R28C34_CE2;
wire R12C6_GB30;
wire R17C32_GB50;
wire R21C23_GB60;
wire R13C3_GB70;
wire R24C24_GBO1;
wire R7C12_GB50;
wire R26C17_GB30;
wire R18C9_GB50;
wire R25C46_GB30;
wire R28C25_N83;
wire R28C43_A6;
wire R22C6_GB40;
wire R6C11_GBO0;
wire R28C40_S80;
wire R26C7_GB50;
wire R24C28_GB60;
wire R7C22_GT10;
wire R5C38_GB40;
wire R11C5_GB00;
wire R14C38_GB70;
wire R24C13_GB60;
wire R3C8_GT00;
wire R6C41_GB30;
wire R10C30_W23;
wire R10C13_E83;
wire R27C29_GBO0;
wire R28C19_X02;
wire R28C31_F5;
wire R5C24_GBO1;
wire R6C38_GT10;
wire R12C21_GB20;
wire R4C7_GB10;
wire R4C17_GB20;
wire R22C2_GB40;
wire R10C16_B4;
wire R29C28_S20;
wire R16C43_GT10;
wire R18C39_GBO0;
wire R10C26_A2;
wire R14C9_GT10;
wire R10C28_SEL1;
wire R2C36_GBO1;
wire R18C8_GB40;
wire R13C10_GB30;
wire R10C10_B7;
wire R28C40_C3;
wire R15C3_GB60;
wire R28C4_CE1;
wire R25C34_GB20;
wire R1C32_E26;
wire R20C2_GB60;
wire R28C43_E21;
wire R5C8_GB50;
wire R10C16_F1;
wire R11C42_GB50;
wire R20C18_SPINE18;
wire R2C22_GT10;
wire R5C37_GBO1;
wire R10C29_N21;
wire R27C17_GBO1;
wire R8C15_GBO1;
wire R2C10_GB70;
wire R6C28_GB30;
wire R12C44_GB70;
wire R10C27_B4;
wire R10C34_W25;
wire R2C15_SPINE9;
wire R9C44_GB20;
wire R14C26_GB50;
wire R14C41_GT10;
wire R7C44_GBO0;
wire R13C8_GB10;
wire R15C25_GB40;
wire R27C23_GB70;
wire R27C44_GB50;
wire R10C29_Q1;
wire R7C18_GB50;
wire R28C34_LSR0;
wire R20C3_SPINE21;
wire R20C37_GBO1;
wire R3C13_GB20;
wire R8C23_GB50;
wire R28C43_B6;
wire R10C26_E10;
wire R14C14_GT00;
wire R18C41_GB60;
wire R27C28_GB50;
wire R10C31_A7;
wire R18C38_GBO1;
wire R4C36_GB10;
wire R16C16_GB60;
wire R16C16_GB00;
wire R28C4_E26;
wire R11C31_GB00;
wire R15C31_GB60;
wire R3C13_GT00;
wire R27C19_GB40;
wire R28C10_W23;
wire R25C8_GB10;
wire R28C7_A1;
wire R28C13_W24;
wire R23C41_GB30;
wire R7C44_GB50;
wire R28C25_W25;
wire R3C22_GBO1;
wire R8C7_GB70;
wire R10C26_Q2;
wire R15C36_GB40;
wire R22C30_GT10;
wire R28C22_N10;
wire R22C40_GB40;
wire R10C37_LSR2;
wire R28C19_C7;
wire R4C42_GBO0;
wire R3C42_GBO1;
wire R2C31_GT00;
wire R6C38_GB10;
wire R1C1_S83;
wire R8C11_GB00;
wire R28C13_C4;
wire R23C34_GB10;
wire R21C2_GB30;
wire R26C37_GBO1;
wire R11C30_GB30;
wire R10C25_E11;
wire R20C14_GB30;
wire R2C30_GB60;
wire R20C29_GB60;
wire R10C28_S13;
wire R12C15_GB70;
wire R28C46_C6;
wire R18C1_GT10;
wire R29C28_SEL2;
wire R29C28_B7;
wire R16C5_GB50;
wire R7C37_GT10;
wire R18C22_GB40;
wire R14C19_GB00;
wire R1C47_A4;
wire R9C17_GBO1;
wire R28C10_A7;
wire R28C13_W27;
wire R6C41_GB00;
wire R26C25_GB60;
wire R1C32_A4;
wire R13C7_GB20;
wire R10C19_X06;
wire R18C29_GB20;
wire R1C47_N25;
wire R17C19_GBO0;
wire R11C23_GT00;
wire R9C5_GB10;
wire R2C18_GB20;
wire R21C14_GB30;
wire R25C14_GB50;
wire R12C23_GB60;
wire R17C43_GB30;
wire R21C11_GB00;
wire R8C42_GB50;
wire R26C29_GB20;
wire R21C35_GB40;
wire R14C33_GB10;
wire R28C4_N26;
wire R11C45_GB00;
wire R28C22_W83;
wire R18C5_GB60;
wire R10C29_N24;
wire R2C37_GBO0;
wire R18C2_GBO1;
wire R5C13_GBO1;
wire R5C26_GB30;
wire R21C23_GB10;
wire R23C40_GB10;
wire R10C27_C4;
wire R26C27_GB50;
wire R8C25_GB40;
wire R14C27_GB10;
wire R26C25_GB10;
wire R1C28_N10;
wire R8C36_GT00;
wire R5C7_GB30;
wire R11C22_GB40;
wire R14C23_GB60;
wire R10C29_S82;
wire R9C5_GT00;
wire R28C22_C7;
wire R7C7_GB50;
wire R5C30_GT00;
wire R18C16_GB10;
wire R17C41_GB00;
wire R18C21_GBO1;
wire R14C31_GB00;
wire R2C43_GB40;
wire R13C19_GB70;
wire R20C31_GB60;
wire R10C10_F0;
wire R10C22_SEL5;
wire R18C9_GB30;
wire R11C27_GB70;
wire R16C37_GBO1;
wire R1C1_D5;
wire R25C42_GT10;
wire R21C35_GT10;
wire R20C17_GB60;
wire R10C27_N12;
wire R15C43_GB30;
wire R15C25_GT10;
wire R10C37_F7;
wire R10C37_F2;
wire R26C27_GB40;
wire R28C4_A2;
wire R16C10_GBO0;
wire R28C37_CLK1;
wire R11C45_GT10;
wire R24C45_GBO1;
wire R18C3_GBO1;
wire R10C19_B7;
wire R15C44_GB10;
wire R23C18_GT10;
wire R10C25_D2;
wire R10C29_X06;
wire R7C40_GBO1;
wire R18C4_GBO1;
wire R3C29_GB50;
wire R21C40_GBO0;
wire R2C35_GT00;
wire R14C31_GT10;
wire R6C18_GT10;
wire R14C2_GB70;
wire R24C4_GB70;
wire R24C24_GB70;
wire R18C31_GB00;
wire R8C20_GB30;
wire R23C22_GB30;
wire R20C32_GB30;
wire R10C40_D3;
wire R22C10_GBO1;
wire R14C17_GT10;
wire R27C37_GBO0;
wire R28C16_CLK1;
wire R8C12_GB20;
wire R4C44_GB30;
wire R10C29_E82;
wire R10C27_F2;
wire R3C40_GBO1;
wire R1C32_E11;
wire R29C28_W83;
wire R4C12_GBO0;
wire R7C18_GB30;
wire R12C27_GB70;
wire R1C47_Q4;
wire R14C41_GB00;
wire R10C40_CLK0;
wire R10C25_SEL4;
wire R20C11_GBO1;
wire R1C28_N82;
wire R10C43_E24;
wire R23C28_GB00;
wire R7C8_GT00;
wire R28C37_B1;
wire R16C17_GB30;
wire R6C27_GB40;
wire R2C32_GB70;
wire R4C26_GB00;
wire R3C6_GB70;
wire R18C2_GT00;
wire R12C38_GB20;
wire R8C43_GT10;
wire R1C1_S11;
wire R17C21_GB70;
wire R11C29_GB00;
wire R22C31_GB00;
wire R12C24_GB10;
wire R5C46_GB20;
wire R10C25_E82;
wire R6C24_GB70;
wire R22C14_GT10;
wire R11C27_GBO0;
wire R10C27_F1;
wire R6C30_GB70;
wire R28C19_N10;
wire R10C10_E80;
wire R12C13_GB40;
wire R17C10_GB70;
wire R6C16_GB50;
wire R16C33_GB00;
wire R20C45_GBO1;
wire R1C47_SEL5;
wire R28C46_B2;
wire R3C21_GB70;
wire R28C13_S81;
wire R28C37_E25;
wire R28C46_SEL7;
wire R9C24_GB70;
wire R6C20_GB40;
wire R10C28_SPINE18;
wire R27C26_GB60;
wire R28C16_SEL1;
wire R28C25_CLK1;
wire R3C20_GB00;
wire R28C40_E80;
wire R26C19_GT00;
wire R3C28_GT10;
wire R5C19_GB50;
wire R13C12_GB40;
wire R16C17_GB70;
wire R14C24_GB60;
wire R7C36_GB70;
wire R25C2_GT10;
wire R17C12_GT10;
wire R10C13_SEL5;
wire R28C22_SEL5;
wire R3C9_GB70;
wire R12C23_GT10;
wire R16C4_GBO1;
wire R12C27_GB00;
wire R23C4_GB40;
wire R12C9_GB20;
wire R18C39_GB60;
wire R24C38_GBO0;
wire R22C33_GB70;
wire R29C28_S12;
wire R18C34_GB20;
wire R20C43_GB10;
wire R16C5_GBO0;
wire R20C11_GB50;
wire R4C21_GB10;
wire R25C16_GB20;
wire R10C30_W13;
wire R21C6_GB00;
wire R24C39_GB10;
wire R28C22_N13;
wire R13C44_GB70;
wire R28C31_N22;
wire R13C22_GB40;
wire R10C27_B2;
wire R18C29_GT10;
wire R1C1_F6;
wire R28C34_Q1;
wire R11C19_GT10;
wire R7C35_GBO1;
wire R7C31_GB70;
wire R14C31_GBO1;
wire R10C25_X04;
wire R10C34_E26;
wire R28C13_N82;
wire R28C7_S21;
wire R7C8_GBO1;
wire R28C4_B2;
wire R10C40_C6;
wire R28C37_C2;
wire R10C34_W20;
wire R13C14_GB60;
wire R9C7_GB60;
wire R9C24_GB60;
wire R10C28_E23;
wire R10C43_Q1;
wire R25C13_GB70;
wire R10C28_S24;
wire R10C43_W81;
wire R10C26_F2;
wire R28C16_E24;
wire R14C7_GBO0;
wire R20C16_GB10;
wire R27C21_GB20;
wire R10C37_N81;
wire R8C21_GBO1;
wire R21C31_GT00;
wire R17C41_GB30;
wire R10C34_SEL5;
wire R20C21_SPINE19;
wire R11C5_GB70;
wire R12C35_GB10;
wire R24C45_GT00;
wire R12C16_GB30;
wire R27C12_GBO1;
wire R2C29_GB50;
wire R17C40_GBO0;
wire R5C19_GB40;
wire R2C35_GB20;
wire R20C37_GB50;
wire R1C28_D5;
wire R28C10_N25;
wire R18C22_GBO0;
wire R16C15_GBO0;
wire R14C8_GBO1;
wire R18C29_GB10;
wire R28C22_E23;
wire R11C29_GB50;
wire R11C11_GB00;
wire R15C6_GB60;
wire R1C32_C5;
wire R13C20_GBO0;
wire R28C28_F4;
wire R4C13_GT00;
wire R14C14_GB30;
wire R4C30_GB20;
wire R13C28_GB00;
wire R8C27_GB70;
wire R10C19_A2;
wire R28C25_E10;
wire R28C16_N81;
wire R11C28_GB30;
wire R21C18_GB20;
wire R14C30_GBO0;
wire R28C13_SEL3;
wire R7C10_GBO0;
wire R23C28_GT00;
wire R18C6_GB00;
wire R5C19_GT00;
wire R9C16_GB20;
wire R24C25_GB50;
wire R23C42_GB60;
wire R10C31_W10;
wire R2C2_GB00;
wire R9C40_GT00;
wire R25C22_GB30;
wire R9C10_GB50;
wire R11C32_GBO1;
wire R20C43_GB60;
wire R15C43_GB70;
wire R18C12_GB50;
wire R28C22_S20;
wire R28C46_S20;
wire R24C17_GBO1;
wire R26C10_GT10;
wire R28C22_B5;
wire R6C13_GB30;
wire R14C27_GB60;
wire R28C46_E27;
wire R11C32_GB10;
wire R9C19_GBO1;
wire R15C9_GB60;
wire R12C46_GB20;
wire R18C11_GB20;
wire R12C28_GB20;
wire R5C30_GB50;
wire R10C26_A6;
wire R28C19_CLK1;
wire R27C8_GB70;
wire R16C31_GB40;
wire R28C4_W24;
wire R1C32_B5;
wire R4C4_GT10;
wire R1C28_D4;
wire R8C7_GB20;
wire R12C24_GB70;
wire R28C4_W26;
wire R28C19_N24;
wire R28C25_CE2;
wire R2C9_SPINE11;
wire R15C32_GB50;
wire R10C29_S11;
wire R25C32_GBO0;
wire R10C30_SPINE1;
wire R20C16_GBO1;
wire R12C12_GB40;
wire R27C35_GT10;
wire R29C28_N10;
wire R10C31_E13;
wire R5C5_GBO0;
wire R10C10_W27;
wire R25C33_GBO0;
wire R6C1_GBO0;
wire R10C27_UNK128;
wire R10C28_W81;
wire R2C19_GBO0;
wire R23C45_GB10;
wire R10C27_W22;
wire R14C34_GBO0;
wire R25C42_GB00;
wire R20C21_GBO1;
wire R10C30_E20;
wire R10C37_F3;
wire R13C40_GB30;
wire R28C25_CE1;
wire R27C44_GT10;
wire R2C2_GB40;
wire R15C7_GB00;
wire R13C32_GB20;
wire R28C34_SEL3;
wire R28C40_F1;
wire R21C8_GB50;
wire R28C22_CLK2;
wire R7C18_GBO1;
wire R28C40_W81;
wire R25C12_GB30;
wire R28C19_W80;
wire R10C29_Q5;
wire R28C22_LSR0;
wire R10C29_A1;
wire R22C5_GB00;
wire R28C16_CE1;
wire R28C34_Q3;
wire R5C25_GB00;
wire R11C25_GB10;
wire R25C20_GB60;
wire R6C32_GB70;
wire R24C15_GB50;
wire R3C19_GB00;
wire R22C3_GB60;
wire R28C46_S11;
wire R27C21_GB40;
wire R16C15_GT10;
wire R8C2_GB20;
wire R26C40_GBO1;
wire R10C29_S25;
wire R8C17_GBO1;
wire R26C1_GBO1;
wire R4C39_GT10;
wire R3C33_GB40;
wire R18C25_GB00;
wire R22C34_GB60;
wire R28C13_E20;
wire R13C6_GT00;
wire R9C24_GB20;
wire R8C19_GB30;
wire R9C31_GB30;
wire R15C7_GB50;
wire R11C14_GB70;
wire R8C37_GBO0;
wire R22C20_GB40;
wire R10C27_F0;
wire R28C4_E23;
wire R27C42_GB20;
wire R10C30_Q3;
wire R22C19_GB40;
wire R3C23_GB40;
wire R18C28_GB20;
wire R27C30_GB40;
wire R16C20_GBO0;
wire R11C19_GB50;
wire R10C16_W20;
wire R10C34_E83;
wire R10C19_B3;
wire R16C36_GB50;
wire R10C30_SEL2;
wire R18C38_GB10;
wire R4C25_GB60;
wire R10C7_E22;
wire R17C36_GB70;
wire R10C13_LSR1;
wire R14C27_GBO0;
wire R10C13_F3;
wire R20C23_GB60;
wire R10C40_S21;
wire R11C41_GB30;
wire R1C1_E24;
wire R16C10_GB00;
wire R10C40_LSR1;
wire R9C39_GB60;
wire R21C44_GB60;
wire R10C28_S23;
wire R28C10_N22;
wire R10C13_X03;
wire R16C28_GB00;
wire R10C29_UNK122;
wire R27C34_GB00;
wire R10C10_E12;
wire R28C10_S82;
wire R4C11_GB20;
wire R8C30_GT00;
wire R17C25_GB10;
wire R12C31_GB30;
wire R22C16_GB40;
wire R5C10_GT10;
wire R8C25_GB10;
wire R10C28_N81;
wire R26C30_GBO1;
wire R2C3_GBO1;
wire R11C41_GT00;
wire R9C41_GB20;
wire R23C27_GBO0;
wire R11C12_GT10;
wire R17C33_GB30;
wire R27C19_GB00;
wire R20C38_GB50;
wire R1C1_Q4;
wire R10C28_C3;
wire R10C34_CE0;
wire R28C34_B3;
wire R25C10_GB30;
wire R28C7_SEL5;
wire R7C25_GBO1;
wire R28C19_W81;
wire R28C40_W24;
wire R24C5_GB00;
wire R24C15_GB20;
wire R17C19_GB30;
wire R14C21_GB60;
wire R3C39_GBO0;
wire R10C26_C0;
wire R23C25_GB70;
wire R16C37_GB30;
wire R7C26_GB00;
wire R7C9_GB10;
wire R25C18_GB10;
wire R16C26_GB10;
wire R20C39_GB20;
wire R6C14_GB30;
wire R13C9_GB10;
wire R18C14_GB60;
wire R22C19_GB60;
wire R17C28_GT10;
wire R4C13_GBO0;
wire R23C20_GB40;
wire R8C20_GBO0;
wire R26C5_GBO0;
wire R17C34_GB00;
wire R16C46_GB20;
wire R20C30_GB40;
wire R23C19_GBO0;
wire R23C31_GBO1;
wire R10C13_A0;
wire R10C19_Q2;
wire R3C9_GBO1;
wire R7C7_GT00;
wire R23C25_GB00;
wire R10C40_Q0;
wire R12C19_GB10;
wire R10C29_S83;
wire R9C7_GB70;
wire R4C32_GT00;
wire R6C12_GBO1;
wire R24C10_GB70;
wire R3C18_GB60;
wire R1C1_X07;
wire R23C42_GB40;
wire R28C7_S80;
wire R22C5_GB50;
wire R1C28_E10;
wire R17C21_GBO0;
wire R27C9_GB60;
wire R2C8_GB40;
wire R14C30_GT00;
wire R18C6_GB10;
wire R10C34_EW10;
wire R5C24_GT00;
wire R11C44_GB70;
wire R21C44_GB50;
wire R5C14_GB30;
wire R18C5_GB50;
wire R17C3_GBO0;
wire R15C9_GB00;
wire R21C28_GB50;
wire R23C43_GB00;
wire R10C31_F0;
wire R18C18_GB40;
wire R23C21_GB40;
wire R5C42_GBO1;
wire R23C28_GB20;
wire R26C19_GB10;
wire R14C29_GB40;
wire R10C28_A5;
wire R28C28_SEL3;
wire R5C11_GB50;
wire R3C33_GBO0;
wire R7C46_GB70;
wire R10C26_S13;
wire R28C40_F7;
wire R29C28_N80;
wire R28C16_W24;
wire R10C29_S81;
wire R3C36_GB30;
wire R11C42_GBO0;
wire R10C30_D4;
wire R28C13_CLK0;
wire R28C28_X08;
wire R5C2_GB20;
wire R28C16_Q4;
wire R28C19_N83;
wire R28C31_S80;
wire R24C25_GB20;
wire R23C20_GB70;
wire R26C21_GB00;
wire R25C38_GB50;
wire R21C41_GB00;
wire R28C40_A6;
wire R28C46_D4;
wire R3C42_GB60;
wire R7C29_GT00;
wire R28C7_S24;
wire R3C26_GB20;
wire R18C13_GT00;
wire R15C44_GT00;
wire R15C40_GB10;
wire R15C44_GBO0;
wire R25C36_GB50;
wire R17C30_GBO1;
wire R9C30_GB30;
wire R10C31_S83;
wire R22C23_GT10;
wire R28C43_S11;
wire R24C29_GB40;
wire R26C7_GB70;
wire R28C7_E20;
wire R28C10_D3;
wire R21C16_GB50;
wire R10C40_B1;
wire R28C16_E26;
wire R28C22_S10;
wire R10C16_B5;
wire R8C33_GBO1;
wire R11C36_GT00;
wire R25C33_GT00;
wire R8C32_GBO1;
wire R16C2_GB60;
wire R18C12_GB70;
wire R23C41_GB10;
wire R24C10_GT00;
wire R20C34_GBO1;
wire R25C24_GB00;
wire R4C34_GB10;
wire R26C26_GB30;
wire R6C41_GB10;
wire R4C3_GBO0;
wire R22C41_GB40;
wire R14C6_GB70;
wire R23C37_GT10;
wire R7C11_GB00;
wire R28C10_W21;
wire R28C19_SN20;
wire R28C7_C4;
wire R24C15_GBO0;
wire R17C15_GT10;
wire R26C11_GBO1;
wire R10C37_C3;
wire R26C35_GB20;
wire R13C12_GB30;
wire R7C18_GT00;
wire R28C34_N82;
wire R16C41_GB60;
wire R28C46_W83;
wire R28C37_W11;
wire R23C8_GB70;
wire R7C4_GB00;
wire R23C21_GT00;
wire R3C6_GBO1;
wire R27C38_GBO0;
wire R10C22_N20;
wire R28C22_E12;
wire R10C26_S80;
wire R28C37_LSR2;
wire R10C16_X07;
wire R17C27_GB50;
wire R25C25_GB70;
wire R10C16_C6;
wire R22C27_GBO1;
wire R2C16_SPINE12;
wire R15C19_GT10;
wire R28C28_N12;
wire R9C44_GT10;
wire R18C30_GB30;
wire R6C42_GBO0;
wire R20C8_GT00;
wire R28C10_SEL4;
wire R28C34_Q6;
wire R11C16_GB60;
wire R9C14_GT10;
wire R10C26_B1;
wire R28C16_E82;
wire R1C47_A0;
wire R25C15_GT00;
wire R11C43_GB30;
wire R22C14_GB00;
wire R4C18_GB50;
wire R11C26_GB70;
wire R22C15_GB10;
wire R5C30_GB20;
wire R21C34_GB10;
wire R18C42_GB10;
wire R21C6_GB60;
wire R28C7_B3;
wire R25C37_GB10;
wire R11C15_GB60;
wire R10C29_D2;
wire R7C23_GB40;
wire R5C34_GB10;
wire R10C27_W80;
wire R1C47_E10;
wire R1C32_X07;
wire R26C44_GT00;
wire R28C25_A6;
wire R18C42_GB70;
wire R2C17_GBO1;
wire R22C33_GB40;
wire R2C37_GB40;
wire R5C6_GB00;
wire R17C11_GT10;
wire R27C12_GB30;
wire R15C26_GBO1;
wire R10C16_CLK0;
wire R26C43_GT10;
wire R23C2_GB00;
wire R12C34_GT00;
wire R18C29_GBO0;
wire R10C40_SEL0;
wire R6C28_GT00;
wire R18C10_GB10;
wire R13C25_GB30;
wire R1C32_Q4;
wire R9C41_GB60;
wire R12C2_GT10;
wire R28C25_S11;
wire R2C2_GB30;
wire R18C44_GT00;
wire R9C9_GB30;
wire R21C34_GB50;
wire R18C20_GB70;
wire R10C28_SEL4;
wire R28C34_E20;
wire R22C7_GB70;
wire R13C22_GB00;
wire R23C13_GB50;
wire R12C40_GB70;
wire R10C19_EW20;
wire R5C17_GT10;
wire R22C44_GBO1;
wire R10C25_W11;
wire R13C28_GB40;
wire R26C32_GBO0;
wire R10C13_D0;
wire R25C46_GB00;
wire R28C22_E83;
wire R16C23_GB70;
wire R22C11_GB30;
wire R28C13_CLK1;
wire R25C17_GB70;
wire R10C27_UNK122;
wire R10C7_Q3;
wire R10C19_S26;
wire R7C26_GB40;
wire R10C34_A6;
wire R22C20_GT00;
wire R28C46_B5;
wire R18C38_GT00;
wire R23C24_GB20;
wire R26C25_GB30;
wire R21C7_GB30;
wire R20C43_GB20;
wire R10C22_SEL3;
wire R20C3_SPINE17;
wire R28C19_S22;
wire R28C31_CLK2;
wire R12C25_GT10;
wire R6C11_GT10;
wire R18C35_GB60;
wire R10C26_E25;
wire R12C19_GB70;
wire R10C37_E20;
wire R24C6_GBO1;
wire R22C43_GBO0;
wire R28C22_W27;
wire R28C40_E21;
wire R5C27_GBO1;
wire R6C2_GBO0;
wire R10C30_C4;
wire R24C9_GB50;
wire R21C36_GB00;
wire R6C26_GB70;
wire R23C29_GB10;
wire R3C28_GT00;
wire R9C22_GB60;
wire R11C26_GB50;
wire R12C20_GT00;
wire R8C34_GB10;
wire R9C42_GB40;
wire R15C40_GBO0;
wire R29C28_A5;
wire R2C20_SPINE12;
wire R28C28_A2;
wire R26C16_GB20;
wire R28C43_N13;
wire R28C7_D1;
wire R27C28_GB00;
wire R24C41_GB40;
wire R2C40_GT10;
wire R3C14_GBO0;
wire R2C17_GB10;
wire R15C8_GT10;
wire R17C15_GB20;
wire R6C35_GB00;
wire R4C10_GB60;
wire R28C19_S24;
wire R1C47_W22;
wire R14C29_GB60;
wire R2C46_GB50;
wire R18C9_GT00;
wire R16C29_GB50;
wire R10C27_D5;
wire R14C37_GB50;
wire R5C3_GB70;
wire R5C9_GB60;
wire R24C19_GBO1;
wire R14C19_GB70;
wire R28C7_S10;
wire R10C7_W22;
wire R12C31_GB50;
wire R1C28_W80;
wire R12C13_GT10;
wire R18C38_GB20;
wire R28C16_E25;
wire R11C7_GBO1;
wire R15C42_GB00;
wire R16C12_GB60;
wire R23C37_GB50;
wire R28C22_B3;
wire R10C13_Q4;
wire R28C13_N24;
wire R10C37_B5;
wire R28C31_W83;
wire R28C25_EW10;
wire R28C37_W23;
wire R12C27_GT10;
wire R5C39_GB00;
wire R26C28_GT00;
wire R5C11_GB70;
wire R16C31_GB70;
wire R10C29_X02;
wire R21C44_GB00;
wire R16C46_GB50;
wire R28C37_D6;
wire R9C23_GB50;
wire R27C29_GB70;
wire R4C27_GB60;
wire R7C2_GB00;
wire R13C8_GB30;
wire R6C25_GB60;
wire R12C7_GB40;
wire R25C8_GB40;
wire R12C5_GB10;
wire R1C28_F0;
wire R22C6_GB20;
wire R21C25_GB30;
wire R10C43_SEL3;
wire R15C26_GB50;
wire R13C35_GBO0;
wire R16C32_GB60;
wire R10C10_Q7;
wire R24C34_GB00;
wire R21C14_GB70;
wire R10C16_B1;
wire R5C5_GB60;
wire R28C13_EW10;
wire R28C34_N80;
wire R1C32_B3;
wire R20C26_GBO0;
wire R28C43_B2;
wire R28C40_E23;
wire R12C33_GBO1;
wire R10C26_SN20;
wire R6C24_GBO1;
wire R6C17_GB50;
wire R7C20_GB10;
wire R20C35_GB50;
wire R27C17_GB60;
wire R15C14_GBO1;
wire R13C7_GB70;
wire R7C46_GB00;
wire R15C6_GBO1;
wire R7C44_GT10;
wire R15C45_GT10;
wire R26C12_GB20;
wire R17C16_GB30;
wire R25C34_GBO0;
wire R22C17_GB10;
wire R15C9_GB40;
wire R21C2_GB10;
wire R17C37_GBO1;
wire R10C19_LSR2;
wire R4C12_GT00;
wire R9C4_GBO0;
wire R10C19_F6;
wire R10C22_S24;
wire R10C27_S11;
wire R14C24_GBO0;
wire R21C37_GBO1;
wire R11C13_GB60;
wire R12C26_GB00;
wire R24C28_GB40;
wire R7C42_GT10;
wire R10C7_Q7;
wire R24C9_GB60;
wire R18C32_GBO0;
wire R13C23_GT10;
wire R10C10_LSR2;
wire R4C20_GB40;
wire R23C44_GB00;
wire R2C12_GB60;
wire R5C21_GB40;
wire R10C13_CE0;
wire R26C9_GB20;
wire R28C19_LSR0;
wire R26C6_GB30;
wire R10C40_S23;
wire R28C10_W12;
wire R11C39_GB40;
wire R4C12_GB70;
wire R13C38_GB10;
wire R27C24_GB40;
wire R20C12_GB00;
wire R16C12_GB30;
wire R12C46_GB70;
wire R14C29_GT00;
wire R25C26_GB30;
wire R14C17_GB40;
wire R13C44_GT00;
wire R25C17_GB40;
wire R10C13_E25;
wire R24C32_GB50;
wire R12C13_GB50;
wire R24C20_GT10;
wire R10C19_CE2;
wire R3C38_GB10;
wire R13C15_GB70;
wire R8C40_GB30;
wire R20C31_GBO0;
wire R28C28_SEL4;
wire R28C37_CE0;
wire R9C18_GB70;
wire R10C28_B2;
wire R20C18_GB70;
wire R10C31_D5;
wire R23C45_GB70;
wire R22C46_GB20;
wire R14C25_GB20;
wire R11C15_GB30;
wire R21C44_GB10;
wire R20C37_SPINE27;
wire R3C13_GT10;
wire R26C13_GB50;
wire R10C27_SEL6;
wire R5C20_GB70;
wire R28C37_W82;
wire R3C10_GB00;
wire R9C40_GB40;
wire R25C30_GBO1;
wire R23C27_GBO1;
wire R6C34_GB40;
wire R22C4_GT10;
wire R8C20_GT10;
wire R21C44_GBO0;
wire R25C8_GBO0;
wire R9C3_GT10;
wire R3C30_GB50;
wire R5C24_GB00;
wire R26C14_GBO0;
wire R21C17_GB50;
wire R10C13_E24;
wire R28C28_X01;
wire R28C43_E82;
wire R8C36_GB50;
wire R22C44_GB00;
wire R10C16_A2;
wire R28C43_N26;
wire R7C24_GB60;
wire R16C12_GB00;
wire R1C28_C5;
wire R15C2_GB20;
wire R10C26_Q1;
wire R27C11_GB40;
wire R16C17_GT10;
wire R20C46_GB10;
wire R27C37_GB00;
wire R20C39_SPINE25;
wire R10C40_X05;
wire R6C20_GBO0;
wire R10C19_F1;
wire R10C43_E81;
wire R24C46_GB50;
wire R10C7_E12;
wire R14C36_GB40;
wire R10C43_S22;
wire R7C4_GB10;
wire R28C10_W22;
wire R10C27_SPINE11;
wire R5C34_GB70;
wire R12C5_GB40;
wire R28C34_W11;
wire R8C23_GB00;
wire R3C29_GT10;
wire R13C4_GB10;
wire R5C45_GB30;
wire R28C4_Q6;
wire R10C7_S27;
wire R28C43_A0;
wire R5C19_GB30;
wire R5C45_GB10;
wire R10C16_N26;
wire R1C32_X05;
wire R21C37_GB10;
wire R15C36_GB20;
wire R28C43_S13;
wire R9C27_GB40;
wire R28C16_S26;
wire R28C25_Q7;
wire R3C12_GBO1;
wire R5C2_GB30;
wire R10C31_Q0;
wire R28C46_C1;
wire R17C35_GB60;
wire R28C13_W25;
wire R15C19_GB30;
wire R29C28_D2;
wire R4C46_GB50;
wire R2C5_GB70;
wire R9C16_GBO0;
wire R4C35_GT00;
wire R3C31_GB00;
wire R16C44_GB40;
wire R2C36_GB30;
wire R21C32_GBO0;
wire R28C31_W81;
wire R9C27_GB50;
wire R11C36_GB00;
wire R24C46_GB60;
wire R25C21_GT10;
wire R28C10_A6;
wire R10C16_C4;
wire R11C3_GT00;
wire R12C12_GB00;
wire R21C24_GB30;
wire R24C35_GT00;
wire R17C21_GB60;
wire R28C10_X06;
wire R5C44_GB10;
wire R25C27_GBO1;
wire R10C13_W22;
wire R12C5_GBO0;
wire R24C22_GB40;
wire R28C13_C3;
wire R14C3_GB00;
wire R14C29_GB20;
wire R9C27_GB30;
wire R27C8_GB50;
wire R23C10_GB60;
wire R23C34_GBO1;
wire R6C31_GB20;
wire R12C40_GB10;
wire R28C31_D4;
wire R12C19_GBO1;
wire R28C25_W82;
wire R28C34_X08;
wire R5C3_GT10;
wire R1C28_E22;
wire R14C36_GBO0;
wire R25C9_GB70;
wire R10C28_X03;
wire R25C2_GB40;
wire R18C12_GBO0;
wire R7C3_GBO1;
wire R13C31_GB50;
wire R29C28_CE2;
wire R24C17_GB30;
wire R2C19_SPINE13;
wire R13C2_GB50;
wire R28C16_X07;
wire R27C10_GB10;
wire R23C29_GB50;
wire R18C22_GB10;
wire R16C31_GB00;
wire R10C31_CLK2;
wire R10C37_N13;
wire R21C9_GB00;
wire R3C17_GBO0;
wire R10C25_Q0;
wire R12C13_GBO1;
wire R16C20_GB40;
wire R28C43_E27;
wire R28C28_W81;
wire R20C7_GT00;
wire R22C3_GB30;
wire R10C43_A0;
wire R28C46_S10;
wire R14C17_GBO0;
wire R12C23_GBO0;
wire R10C7_X04;
wire R26C24_GB30;
wire R14C31_GB30;
wire R28C13_E11;
wire R7C6_GT10;
wire R12C25_GB50;
wire R23C15_GT10;
wire R27C34_GB50;
wire R28C22_W22;
wire R27C36_GBO0;
wire R28C22_EW10;
wire R28C25_W10;
wire R27C45_GB70;
wire R9C25_GB20;
wire R10C30_N10;
wire R10C30_S13;
wire R26C29_GB40;
wire R13C6_GB30;
wire R10C22_A0;
wire R11C29_GT10;
wire R11C45_GB70;
wire R6C3_GB30;
wire R10C34_B1;
wire R11C24_GB20;
wire R28C28_X06;
wire R17C36_GB00;
wire R23C38_GB20;
wire R8C32_GT10;
wire R20C17_GB10;
wire R10C7_E23;
wire R10C27_F4;
wire R28C31_W11;
wire R17C45_GB40;
wire R14C23_GB20;
wire R22C7_GBO0;
wire R4C40_GB20;
wire R10C7_D1;
wire R28C43_W83;
wire R10C26_B0;
wire R10C27_W25;
wire R28C46_S83;
wire R28C4_Q4;
wire R28C4_N83;
wire R15C32_GB00;
wire R16C17_GT00;
wire R1C1_E10;
wire R3C4_GB30;
wire R5C12_GBO1;
wire R18C16_GB40;
wire R4C16_GB30;
wire R24C17_GB70;
wire R25C25_GT10;
wire R10C28_F0;
wire R18C6_GB40;
wire R18C23_GB20;
wire R25C40_GB50;
wire R28C19_B2;
wire R23C1_GT00;
wire R1C1_N23;
wire R10C25_S27;
wire R15C1_GT10;
wire R21C28_GB10;
wire R12C6_GB20;
wire R24C25_GB60;
wire R4C12_GB20;
wire R6C38_GBO1;
wire R4C8_GBO1;
wire R24C5_GT10;
wire R26C38_GBO0;
wire R10C28_N20;
wire R10C31_N25;
wire R16C37_GT10;
wire R2C36_GB10;
wire R4C10_GB50;
wire R15C26_GB00;
wire R28C19_E27;
wire R17C5_GB60;
wire R27C41_GB10;
wire R11C39_GB20;
wire R27C4_GB50;
wire R23C7_GB20;
wire R25C35_GT10;
wire R16C33_GB70;
wire R22C16_GT10;
wire R10C29_W12;
wire R28C31_W27;
wire R17C5_GT10;
wire R10C7_C1;
wire R26C22_GB40;
wire R10C22_B0;
wire R5C22_GT00;
wire R10C27_S21;
wire R18C10_GB70;
wire R10C43_LSR1;
wire R22C26_GB70;
wire R10C25_S23;
wire R10C19_E21;
wire R20C27_GB70;
wire R27C34_GT10;
wire R8C9_GBO0;
wire R26C8_GT10;
wire R8C3_GB50;
wire R23C24_GB40;
wire R10C34_CLK2;
wire R28C4_S81;
wire R2C15_GB30;
wire R2C3_GB30;
wire R24C15_GB00;
wire R28C43_E24;
wire R7C17_GB70;
wire R29C28_S11;
wire R8C3_GB10;
wire R16C23_GB50;
wire R17C44_GB60;
wire R4C6_GT00;
wire R28C46_D0;
wire R22C40_GBO1;
wire R8C15_GB50;
wire R26C32_GB10;
wire R10C27_X06;
wire R21C26_GB00;
wire R17C40_GB70;
wire R25C46_GB20;
wire R7C16_GB10;
wire R13C33_GB10;
wire R25C36_GB70;
wire R27C44_GB60;
wire R28C7_E21;
wire R3C23_GB60;
wire R14C46_GT00;
wire R27C28_GB60;
wire R11C38_GB40;
wire R10C43_X04;
wire R24C7_GBO1;
wire R8C41_GB20;
wire R10C13_N80;
wire R25C25_GT00;
wire R22C45_GT00;
wire R11C30_GB20;
wire R5C32_GB30;
wire R6C6_GB10;
wire R28C34_E27;
wire R10C22_S83;
wire R18C34_GB00;
wire R28C4_W20;
wire R20C15_GBO1;
wire R9C29_GB00;
wire R28C46_N11;
wire R20C32_GB40;
wire R25C3_GB20;
wire R23C7_GB40;
wire R26C39_GB30;
wire R2C40_SPINE0;
wire R11C18_GB60;
wire R10C26_Q7;
wire R16C22_GB20;
wire R24C13_GT00;
wire R26C19_GT10;
wire R24C32_GT00;
wire R4C17_GBO0;
wire R12C20_GB70;
wire R11C26_GB10;
wire R20C9_SPINE19;
wire R11C31_GT00;
wire R18C42_GT00;
wire R21C16_GB20;
wire R2C19_GB50;
wire R11C40_GB10;
wire R10C34_SN20;
wire R26C17_GB20;
wire R13C20_GT10;
wire R3C39_GB50;
wire R28C46_N80;
wire R22C18_GT00;
wire R20C29_GB20;
wire R20C39_GB70;
wire R10C13_S25;
wire R28C7_A0;
wire R2C19_GB30;
wire R20C36_GB00;
wire R10C30_N21;
wire R6C33_GB00;
wire R6C2_GB50;
wire R25C10_GB50;
wire R28C22_E80;
wire R24C21_GT00;
wire R4C6_GB20;
wire R7C40_GT10;
wire R7C21_GBO0;
wire R5C13_GB30;
wire R2C15_GB20;
wire R10C10_N23;
wire R21C33_GB00;
wire R10C10_N26;
wire R13C27_GB50;
wire R3C38_GB20;
wire R22C29_GB20;
wire R10C10_F3;
wire R8C13_GB40;
wire R9C23_GB30;
wire R13C16_GB00;
wire R3C12_GB40;
wire R20C15_GB70;
wire R13C46_GB10;
wire R10C28_S82;
wire R11C43_GT00;
wire R28C10_C2;
wire R27C6_GB20;
wire R10C10_X08;
wire R15C35_GT00;
wire R6C19_GB50;
wire R5C34_GBO0;
wire R11C42_GB30;
wire R3C20_GT10;
wire R24C16_GB40;
wire R15C34_GB10;
wire R4C22_GB40;
wire R5C36_GT10;
wire R17C38_GB70;
wire R10C31_X01;
wire R1C28_EW10;
wire R28C19_S13;
wire R26C9_GB00;
wire R17C26_GBO1;
wire R3C19_GB50;
wire R9C27_GB10;
wire R10C34_LSR2;
wire R2C38_GT10;
wire R2C2_GBO1;
wire R21C19_GB20;
wire R20C19_SPINE17;
wire R22C26_GB40;
wire R4C31_GBO0;
wire R9C5_GB40;
wire R3C30_GBO0;
wire R17C13_GBO1;
wire R24C32_GB10;
wire R21C2_GB60;
wire R23C36_GB10;
wire R12C40_GB60;
wire R22C10_GB40;
wire R10C19_W22;
wire R26C6_GB10;
wire R1C32_N81;
wire R10C19_Q6;
wire R10C29_B1;
wire R11C38_GT00;
wire R18C18_GB20;
wire R27C29_GB40;
wire R27C37_GB20;
wire R23C11_GT10;
wire R18C5_GB70;
wire R12C30_GBO1;
wire R23C22_GB10;
wire R5C19_GB20;
wire R26C14_GB70;
wire R20C39_GB50;
wire R6C16_GT00;
wire R22C12_GBO1;
wire R10C7_E10;
wire R10C29_F7;
wire R6C17_GT00;
wire R10C30_LSR0;
wire R21C28_GB20;
wire R27C27_GB30;
wire R4C43_GBO1;
wire R10C29_S20;
wire R10C40_W22;
wire R28C34_N25;
wire R20C7_GB10;
wire R1C1_S82;
wire R27C34_GB40;
wire R1C32_N24;
wire R27C20_GB30;
wire R1C47_D0;
wire R10C37_CE1;
wire R23C21_GB60;
wire R21C38_GT00;
wire R26C18_GB70;
wire R15C9_GB30;
wire R4C31_GB10;
wire R28C25_SEL2;
wire R28C22_E13;
wire R15C44_GB60;
wire R28C4_N23;
wire R1C32_Q7;
wire R10C30_E12;
wire R10C29_S13;
wire R28C40_N20;
wire R6C23_GB10;
wire R24C13_GB20;
wire R12C12_GB70;
wire R10C26_SEL0;
wire R18C16_GT00;
wire R2C45_GBO1;
wire R20C27_GB20;
wire R8C32_GB10;
wire R28C37_W26;
wire R14C24_GB00;
wire R7C3_GT10;
wire R28C13_D6;
wire R10C16_N82;
wire R10C28_E25;
wire R24C39_GBO0;
wire R14C16_GB50;
wire R22C9_GB50;
wire R2C12_GB30;
wire R4C3_GB50;
wire R28C4_N13;
wire R20C4_GT10;
wire R21C39_GT10;
wire R9C40_GBO0;
wire R12C30_GB50;
wire R18C1_GBO0;
wire R4C27_GBO1;
wire R18C25_GB20;
wire R13C9_GB70;
wire R13C35_GB20;
wire R28C7_C1;
wire R10C19_Q5;
wire R10C43_E12;
wire R6C22_GB40;
wire R10C28_A3;
wire R18C23_GB40;
wire R4C30_GB70;
wire R10C28_W80;
wire R1C47_E80;
wire R11C3_GB70;
wire R26C30_GB00;
wire R10C25_CE2;
wire R10C27_S83;
wire R17C47_F6;
wire R18C35_GB50;
wire R4C14_GB60;
wire R10C26_SEL6;
wire R5C7_GT10;
wire R5C12_GB20;
wire R25C7_GBO0;
wire R16C3_GB20;
wire R22C39_GB70;
wire R24C31_GB60;
wire R10C10_C2;
wire R10C22_C6;
wire R28C19_SEL4;
wire R10C30_D0;
wire R15C2_GT10;
wire R28C13_SEL6;
wire R5C38_GB20;
wire R20C6_GB50;
wire R2C29_GB00;
wire R25C22_GBO1;
wire R22C13_GB60;
wire R15C15_GB70;
wire R25C7_GB20;
wire R22C18_GB20;
wire R29C28_E23;
wire R28C31_C2;
wire R27C6_GB50;
wire R1C32_W81;
wire R3C21_GB60;
wire R15C38_GB00;
wire R26C13_GB20;
wire R13C32_GT10;
wire R26C16_GB70;
wire R22C31_GBO0;
wire R11C46_GBO0;
wire R10C34_SEL1;
wire R2C8_GT10;
wire R29C28_D7;
wire R24C42_GBO1;
wire R13C45_GBO1;
wire R13C38_GB20;
wire R27C3_GT10;
wire R28C25_S21;
wire R6C11_GB40;
wire R3C27_GB10;
wire R14C17_GB20;
wire R16C27_GB20;
wire R5C4_GB10;
wire R26C9_GBO0;
wire R26C20_GB50;
wire R28C25_F4;
wire R14C8_GT10;
wire R13C8_GBO1;
wire R23C39_GB20;
wire R21C25_GB50;
wire R8C11_GB50;
wire R22C46_GBO1;
wire R10C16_E25;
wire R17C43_GT00;
wire R27C15_GB20;
wire R28C25_C5;
wire R9C22_GBO0;
wire R20C4_GB50;
wire R26C38_GB50;
wire R25C16_GB00;
wire R18C23_GB10;
wire R7C41_GB50;
wire R16C43_GB10;
wire R10C22_E27;
wire R6C3_GB60;
wire R25C37_GB20;
wire R10C34_B6;
wire R28C19_CLK2;
wire R28C34_SN10;
wire R2C8_GB30;
wire R12C41_GT10;
wire R9C16_GB40;
wire R26C20_GT10;
wire R1C28_A1;
wire R4C23_GB60;
wire R10C19_S22;
wire R6C3_GBO1;
wire R22C27_GB20;
wire R11C39_GB70;
wire R25C42_GB60;
wire R10C22_F0;
wire R10C31_F2;
wire R28C7_E25;
wire R16C44_GB00;
wire R9C42_GBO0;
wire R28C13_X07;
wire R26C43_GT00;
wire R6C16_GB40;
wire R24C30_GB10;
wire R12C25_GT00;
wire R4C45_GBO1;
wire R15C10_GBO0;
wire R7C38_GBO1;
wire R2C24_GBO1;
wire R14C2_GB00;
wire R26C36_GB60;
wire R17C16_GB10;
wire R13C38_GBO0;
wire R23C31_GB00;
wire R28C16_C0;
wire R16C37_GB10;
wire R2C38_SPINE2;
wire R7C26_GT00;
wire R21C23_GB30;
wire R18C17_GB70;
wire R4C39_GB00;
wire R11C19_GT00;
wire R13C13_GB50;
wire R6C45_GB00;
wire R20C2_GB50;
wire R10C25_SEL2;
wire R28C28_B2;
wire R20C20_GB00;
wire R21C20_GB10;
wire R12C10_GB60;
wire R8C19_GB20;
wire R3C28_GB40;
wire R15C41_GB60;
wire R26C9_GB30;
wire R10C10_E26;
wire R25C15_GT10;
wire R10C26_W22;
wire R25C12_GT10;
wire R5C8_GB60;
wire R7C21_GB30;
wire R28C31_N25;
wire R3C9_GB20;
wire R8C9_GT00;
wire R13C43_GB70;
wire R5C8_GBO1;
wire R22C40_GB10;
wire R10C7_N81;
wire R18C16_GT10;
wire R3C8_GB50;
wire R16C9_GB00;
wire R13C20_GB30;
wire R13C6_GB40;
wire R28C37_A1;
wire R5C13_GBO0;
wire R5C44_GB30;
wire R20C34_GB20;
wire R20C29_SPINE27;
wire R25C44_GBO0;
wire R4C15_GBO1;
wire R25C3_GB00;
wire R23C10_GB10;
wire R28C34_S20;
wire R22C14_GB20;
wire R11C17_GT10;
wire R10C7_S12;
wire R11C11_GT00;
wire R2C16_GBO0;
wire R9C26_GT10;
wire R3C20_GB50;
wire R22C27_GB50;
wire R16C41_GT00;
wire R28C4_E10;
wire R5C36_GBO0;
wire R28C31_Q1;
wire R28C16_N80;
wire R28C28_Q2;
wire R17C43_GB10;
wire R4C16_GB20;
wire R13C4_GBO1;
wire R28C7_Q3;
wire R3C41_GBO0;
wire R28C43_CLK1;
wire R20C6_GB00;
wire R5C29_GB40;
wire R27C36_GB30;
wire R6C30_GB30;
wire R10C28_D7;
wire R10C22_EW20;
wire R24C38_GB60;
wire R22C38_GT00;
wire R14C11_GBO0;
wire R13C5_GBO0;
wire R10C19_S82;
wire R25C5_GB30;
wire R9C35_GB00;
wire R18C25_GBO0;
wire R13C38_GB30;
wire R21C27_GB20;
wire R10C13_E23;
wire R28C34_N27;
wire R16C25_GT00;
wire R28C22_Q0;
wire R1C32_N22;
wire R12C31_GBO0;
wire R13C27_GB30;
wire R10C37_SN10;
wire R28C22_N24;
wire R28C31_F7;
wire R10C7_X05;
wire R20C21_GB50;
wire R17C10_GT00;
wire R10C34_X02;
wire R29C28_E26;
wire R9C13_GT10;
wire R21C17_GB40;
wire R13C37_GBO0;
wire R12C39_GBO1;
wire R14C41_GBO1;
wire R15C26_GT00;
wire R14C8_GB60;
wire R10C34_D0;
wire R7C37_GB40;
wire R28C31_X05;
wire R21C13_GT00;
wire R28C4_SEL4;
wire R8C13_GB60;
wire R23C29_GB40;
wire R28C28_N23;
wire R10C10_W26;
wire R12C20_GB10;
wire R28C22_E27;
wire R1C32_E12;
wire R10C10_B0;
wire R10C28_N82;
wire R10C40_W80;
wire R10C31_E20;
wire R28C4_N81;
wire R23C13_GBO0;
wire R28C34_SEL5;
wire R18C15_GB50;
wire R21C30_GB40;
wire R18C4_GB00;
wire R10C13_B6;
wire R1C47_N26;
wire R14C18_GBO0;
wire R8C46_GB50;
wire R3C1_GT10;
wire R13C26_GT00;
wire R12C19_GB20;
wire R24C40_GB40;
wire R10C19_N11;
wire R28C4_S80;
wire R2C21_GB60;
wire R4C45_GB10;
wire R8C24_GB40;
wire R18C23_GB50;
wire R10C27_Q6;
wire R21C27_GB50;
wire R17C23_GB70;
wire R3C4_GT10;
wire R13C3_GB10;
wire R15C1_GBO0;
wire R24C14_GB70;
wire R9C38_GT00;
wire R11C46_GB00;
wire R24C44_GB30;
wire R27C4_GB00;
wire R7C38_GB30;
wire R23C39_GB50;
wire R10C13_SEL7;
wire R14C43_GB50;
wire R25C26_GB70;
wire R27C35_GB20;
wire R4C45_GT00;
wire R17C10_GB30;
wire R10C31_A3;
wire R17C18_GT10;
wire R23C2_GB10;
wire R6C36_GB00;
wire R8C36_GB30;
wire R10C43_S21;
wire R28C4_CLK1;
wire R2C32_GBO1;
wire R1C28_W25;
wire R24C9_GT10;
wire R10C34_X04;
wire R16C20_GB20;
wire R9C4_GB00;
wire R22C2_GB60;
wire R10C27_C6;
wire R10C22_W24;
wire R2C37_GB60;
wire R1C28_SEL0;
wire R1C28_D7;
wire R27C23_GT10;
wire R6C16_GB70;
wire R15C26_GT10;
wire R2C7_GT00;
wire R24C22_GT10;
wire R11C36_GB70;
wire R28C7_N26;
wire R27C25_GT10;
wire R15C8_GBO0;
wire R10C34_E82;
wire R18C15_GB30;
wire R15C23_GT10;
wire R17C22_GB00;
wire R10C34_S81;
wire R8C21_GB40;
wire R14C20_GB10;
wire R8C40_GT00;
wire R13C6_GB00;
wire R16C40_GB70;
wire R3C46_GB40;
wire R10C30_N83;
wire R10C40_SEL4;
wire R15C17_GT10;
wire R10C30_A5;
wire R16C7_GB30;
wire R28C25_C2;
wire R17C8_GB40;
wire R20C16_SPINE20;
wire R24C27_GB20;
wire R18C20_GB40;
wire R27C35_GB50;
wire R27C33_GB30;
wire R21C8_GT00;
wire R24C39_GB00;
wire R24C42_GB10;
wire R9C23_GB70;
wire R2C35_GB70;
wire R7C38_GBO0;
wire R28C4_SEL3;
wire R26C39_GB00;
wire R7C19_GT00;
wire R18C39_GB20;
wire R9C22_GB10;
wire R15C14_GBO0;
wire R8C6_GB70;
wire R3C20_GT00;
wire R8C9_GB70;
wire R15C28_GB30;
wire R23C14_GB40;
wire R11C2_GBO1;
wire R25C22_GB00;
wire R10C31_W25;
wire R7C9_GB70;
wire R4C37_GB00;
wire R10C40_A3;
wire R20C15_SPINE17;
wire R9C10_GB30;
wire R28C4_F4;
wire R25C6_GB50;
wire R9C14_GB10;
wire R2C25_GB70;
wire R24C25_GB30;
wire R10C22_D5;
wire R6C31_GB10;
wire R10C29_E21;
wire R12C41_GB00;
wire R4C21_GT00;
wire R22C42_GBO1;
wire R5C42_GB50;
wire R27C16_GB40;
wire R4C16_GT10;
wire R27C29_GB00;
wire R28C46_N10;
wire R13C31_GB30;
wire R1C28_D3;
wire R27C46_GB60;
wire R28C46_E10;
wire R18C43_GB10;
wire R28C28_C0;
wire R25C40_GB60;
wire R25C21_GB00;
wire R8C26_GB20;
wire R11C29_GBO1;
wire R3C36_GBO1;
wire R5C36_GB50;
wire R23C31_GBO0;
wire R2C31_SPINE5;
wire R9C26_GB60;
wire R1C1_F5;
wire R16C45_GBO1;
wire R6C24_GB10;
wire R28C28_W26;
wire R24C39_GB30;
wire R10C7_SEL2;
wire R22C45_GB60;
wire R23C8_GBO0;
wire R10C30_SEL0;
wire R8C33_GB30;
wire R28C13_SEL4;
wire R8C34_GB70;
wire R22C7_GB50;
wire R22C15_GB40;
wire R8C38_GB50;
wire R10C22_S12;
wire R28C13_A1;
wire R10C31_S10;
wire R10C13_S83;
wire R10C28_S21;
wire R11C6_GB30;
wire R17C4_GBO0;
wire R25C38_GB70;
wire R1C47_E12;
wire R17C39_GB10;
wire R1C28_W21;
wire R29C28_SN20;
wire R1C47_W25;
wire R1C28_W10;
wire R1C32_LSR1;
wire R10C7_A5;
wire R20C40_SPINE28;
wire R7C17_GBO0;
wire R9C6_GT00;
wire R26C31_GB70;
wire R7C32_GBO1;
wire R3C6_GT10;
wire R24C8_GB30;
wire R15C3_GT10;
wire R25C12_GB70;
wire R15C25_GB20;
wire R9C30_GB70;
wire R15C23_GT00;
wire R14C2_GB50;
wire R21C38_GB70;
wire R21C39_GB50;
wire R11C6_GT00;
wire R27C14_GBO0;
wire R10C28_SEL3;
wire R10C34_C2;
wire R15C15_GBO1;
wire R12C2_GB60;
wire R10C40_A7;
wire R28C16_S82;
wire R16C19_GBO0;
wire R15C7_GB40;
wire R10C25_A7;
wire R28C19_N21;
wire R29C28_A3;
wire R4C10_GT00;
wire R6C21_GBO0;
wire R4C26_GB70;
wire R28C16_X03;
wire R17C37_GB40;
wire R4C24_GB50;
wire R7C41_GB60;
wire R4C42_GB70;
wire R27C46_GB40;
wire R28C43_E10;
wire R26C10_GB40;
wire R28C7_N21;
wire R21C42_GB40;
wire R7C41_GB40;
wire R10C30_B7;
wire R13C34_GB40;
wire R8C36_GB40;
wire R28C34_W12;
wire R10C31_F5;
wire R7C13_GB70;
wire R13C44_GB30;
wire R26C35_GT00;
wire R17C4_GB40;
wire R7C32_GB10;
wire R28C46_Q5;
wire R11C26_GB20;
wire R6C24_GB40;
wire R17C10_GBO0;
wire R17C40_GB20;
wire R16C27_GT00;
wire R28C46_E83;
wire R10C40_C7;
wire R1C28_W24;
wire R10C19_E10;
wire R8C27_GB00;
wire R5C18_GT10;
wire R21C45_GB70;
wire R9C24_GT10;
wire R28C46_C7;
wire R13C30_GBO0;
wire R10C29_B3;
wire R22C24_GBO0;
wire R10C25_Q7;
wire R17C2_GB00;
wire R18C32_GB10;
wire R6C6_GBO1;
wire R26C44_GB00;
wire R1C1_W10;
wire R3C7_GB20;
wire R10C19_C4;
wire R20C11_GB20;
wire R27C11_GB00;
wire R8C11_GBO1;
wire R26C33_GB70;
wire R2C10_GB10;
wire R23C14_GB50;
wire R10C37_Q3;
wire R22C10_GB10;
wire R11C6_GBO0;
wire R28C22_W23;
wire R23C7_GT10;
wire R23C24_GB30;
wire R10C27_S12;
wire R17C20_GB50;
wire R14C32_GB10;
wire R12C41_GB20;
wire R16C17_GB10;
wire R12C27_GBO0;
wire R22C24_GB60;
wire R15C42_GB30;
wire R14C12_GB70;
wire R10C7_CLK0;
wire R10C26_W20;
wire R28C16_W21;
wire R10C25_D7;
wire R28C19_SEL7;
wire R22C13_GBO1;
wire R7C4_GB30;
wire R20C20_GB60;
wire R10C7_N23;
wire R24C32_GB00;
wire R15C11_GB00;
wire R28C7_A2;
wire R28C10_W25;
wire R28C37_W22;
wire R26C8_GB50;
wire R29C28_W20;
wire R18C16_GBO1;
wire R15C41_GB00;
wire R24C34_GBO1;
wire R10C22_D0;
wire R20C34_GB70;
wire R20C24_GB60;
wire R28C34_D6;
wire R10C13_EW20;
wire R11C34_GB20;
wire R7C39_GT00;
wire R13C19_GT10;
wire R29C28_F2;
wire R22C22_GBO0;
wire R6C12_GB60;
wire R14C28_GT00;
wire R10C22_E82;
wire R9C39_GB10;
wire R8C1_GBO0;
wire R7C9_GBO1;
wire R18C2_GBO0;
wire R17C24_GB50;
wire R10C28_A6;
wire R28C25_N26;
wire R10C31_SN20;
wire R17C40_GT00;
wire R16C9_GBO0;
wire R26C5_GB20;
wire R28C46_W23;
wire R5C7_GB50;
wire R9C27_GBO0;
wire R29C28_CE1;
wire R8C23_GB20;
wire R27C27_GBO0;
wire R25C13_GB60;
wire R26C36_GB70;
wire R28C34_B5;
wire R12C2_GT00;
wire R5C31_GBO1;
wire R9C32_GB50;
wire R25C41_GB50;
wire R28C37_W27;
wire R23C14_GB70;
wire R20C13_GB30;
wire R15C42_GB10;
wire R21C2_GBO0;
wire R1C1_A0;
wire R10C37_SEL1;
wire R8C30_GB50;
wire R10C37_E81;
wire R26C30_GT00;
wire R15C19_GB50;
wire R6C35_GBO1;
wire R21C22_GBO0;
wire R20C5_GT00;
wire R3C7_GB30;
wire R20C45_GB40;
wire R24C33_GBO1;
wire R1C32_SEL6;
wire R29C28_E12;
wire R1C47_E83;
wire R7C27_GBO1;
wire R21C10_GT10;
wire R21C41_GB10;
wire R17C8_GBO0;
wire R8C41_GB40;
wire R10C30_SN10;
wire R3C36_GB60;
wire R28C46_B1;
wire R7C25_GB40;
wire R28C28_W83;
wire R26C33_GB30;
wire R9C14_GB40;
wire R13C45_GB40;
wire R3C6_GB60;
wire R10C16_SEL4;
wire R10C25_B6;
wire R15C40_GBO1;
wire R2C20_GT00;
wire R2C5_GBO0;
wire R4C9_GB70;
wire R20C10_GB60;
wire R3C46_GB10;
wire R3C37_GB60;
wire R18C41_GB10;
wire R12C35_GB70;
wire R10C28_D6;
wire R3C43_GB60;
wire R24C6_GB00;
wire R15C21_GB30;
wire R28C40_EW10;
wire R9C42_GB60;
wire R20C39_GB00;
wire R14C39_GBO1;
wire R8C27_GB30;
wire R12C44_GB30;
wire R28C34_Q2;
wire R28C16_SEL0;
wire R25C41_GB20;
wire R11C16_GB10;
wire R20C31_GB40;
wire R16C28_GB10;
wire R23C9_GT00;
wire R10C30_W80;
wire R28C34_CE0;
wire R20C8_GB30;
wire R9C17_GB10;
wire R18C32_GB30;
wire R16C6_GB60;
wire R8C25_GB20;
wire R17C19_GT10;
wire R9C9_GB60;
wire R10C30_S26;
wire R5C24_GB60;
wire R22C27_GB70;
wire R26C6_GB50;
wire R28C4_A5;
wire R28C43_LSR2;
wire R5C3_GB40;
wire R11C43_GB40;
wire R10C25_W27;
wire R3C3_GB10;
wire R28C4_CE0;
wire R16C3_GB00;
wire R20C10_GT10;
wire R28C25_W80;
wire R10C7_E81;
wire R22C10_GT10;
wire R4C19_GB20;
wire R28C40_Q2;
wire R10C28_CE1;
wire R3C17_GB20;
wire R16C18_GB50;
wire R1C28_W11;
wire R14C15_GB40;
wire R10C10_F6;
wire R5C15_GBO0;
wire R28C46_E81;
wire R5C12_GB50;
wire R1C28_CLK2;
wire R10C22_E26;
wire R21C42_GB60;
wire R24C19_GB60;
wire R11C6_GBO1;
wire R24C40_GT10;
wire R16C24_GB00;
wire R10C27_S80;
wire R2C22_GB50;
wire R10C43_B0;
wire R28C19_SN10;
wire R17C17_GB30;
wire R27C21_GBO1;
wire R24C19_GB70;
wire R1C1_N25;
wire R8C17_GB20;
wire R23C44_GT10;
wire R24C35_GB20;
wire R11C31_GB50;
wire R6C29_GB30;
wire R27C42_GB50;
wire R13C37_GT10;
wire R20C2_GB00;
wire R27C34_GBO0;
wire R18C44_GB20;
wire R26C3_GBO0;
wire R10C26_E27;
wire R5C46_GB50;
wire R16C35_GB00;
wire R28C22_CLK1;
wire R24C46_GBO1;
wire R10C26_C4;
wire R8C41_GB30;
wire R8C45_GB40;
wire R14C34_GB30;
wire R13C11_GB70;
wire R8C6_GB10;
wire R17C16_GB20;
wire R24C21_GB40;
wire R22C20_GBO0;
wire R15C23_GBO0;
wire R7C1_GBO1;
wire R12C18_GB30;
wire R10C26_SEL7;
wire R16C27_GBO0;
wire R24C6_GBO0;
wire R10C25_N10;
wire R8C29_GB70;
wire R18C2_GB30;
wire R28C43_X03;
wire R21C16_GT10;
wire R14C7_GB40;
wire R3C21_GBO0;
wire R16C30_GB40;
wire R20C28_GB00;
wire R11C36_GBO1;
wire R10C10_W23;
wire R21C37_GB30;
wire R28C43_W20;
wire R28C25_C3;
wire R9C13_GBO1;
wire R18C40_GB20;
wire R3C16_GB60;
wire R21C19_GB30;
wire R21C25_GB60;
wire R10C26_LSR2;
wire R21C37_GB70;
wire R10C13_W23;
wire R25C4_GB30;
wire R3C40_GB10;
wire R2C29_GB10;
wire R15C14_GB60;
wire R7C37_GB00;
wire R2C29_GBO0;
wire R10C7_A1;
wire R9C25_GT00;
wire R16C20_GB30;
wire R26C31_GB10;
wire R28C22_F6;
wire R8C40_GB70;
wire R12C36_GBO0;
wire R10C13_N26;
wire R5C13_GB60;
wire R2C30_GB00;
wire R17C36_GB30;
wire R23C11_GB10;
wire R22C12_GT10;
wire R10C27_SN10;
wire R17C2_GB30;
wire R18C35_GB30;
wire R15C5_GBO1;
wire R28C40_SEL2;
wire R10C7_N27;
wire R18C34_GB40;
wire R17C18_GB70;
wire R1C28_A6;
wire R12C39_GBO0;
wire R23C35_GB10;
wire R10C43_W83;
wire R22C26_GB30;
wire R1C32_N20;
wire R20C17_SPINE19;
wire R27C27_GB20;
wire R16C13_GBO0;
wire R26C14_GBO1;
wire R14C37_GB40;
wire R5C14_GB70;
wire R21C19_GB60;
wire R22C33_GB10;
wire R3C29_GB00;
wire R20C20_SPINE16;
wire R25C18_GT00;
wire R14C21_GB50;
wire R10C37_C2;
wire R18C23_GB30;
wire R15C13_GT00;
wire R10C30_A2;
wire R7C30_GB40;
wire R13C46_GB40;
wire R10C22_X05;
wire R2C9_GBO1;
wire R4C40_GB40;
wire R23C31_GB10;
wire R27C22_GBO1;
wire R17C6_GB30;
wire R23C3_GT00;
wire R23C8_GB50;
wire R7C44_GT00;
wire R13C38_GB50;
wire R12C2_GBO0;
wire R20C14_GB60;
wire R28C4_W21;
wire R27C24_GT10;
wire R24C10_GBO0;
wire R10C16_CLK2;
wire R1C1_E80;
wire R8C28_GT10;
wire R13C4_GB20;
wire R10C29_S27;
wire R27C21_GB50;
wire R6C37_GT00;
wire R28C37_SEL1;
wire R8C26_GBO1;
wire R11C35_GT00;
wire R29C28_S26;
wire R1C1_W25;
wire R27C13_GB10;
wire R23C45_GBO1;
wire R28C7_E12;
wire R3C29_GB70;
wire R3C25_GB30;
wire R15C8_GB70;
wire R10C25_C1;
wire R14C16_GB00;
wire R10C28_F3;
wire R25C13_GB50;
wire R28C22_F1;
wire R4C4_GBO1;
wire R28C10_A4;
wire R28C25_X05;
wire R4C38_GB70;
wire R27C15_GT00;
wire R14C41_GB30;
wire R27C45_GB40;
wire R28C37_F3;
wire R2C32_GB20;
wire R10C34_E81;
wire R28C7_W82;
wire R10C34_X05;
wire R17C40_GB50;
wire R3C43_GB20;
wire R27C34_GT00;
wire R5C6_GB20;
wire R26C24_GB50;
wire R25C21_GBO1;
wire R8C41_GB60;
wire R4C44_GB40;
wire R28C34_S10;
wire R10C13_C7;
wire R3C2_GB40;
wire R4C20_GBO1;
wire R12C34_GB10;
wire R3C17_GT10;
wire R28C7_C6;
wire R7C30_GB30;
wire R2C33_GB60;
wire R22C6_GT00;
wire R13C23_GBO1;
wire R2C4_GBO0;
wire R7C6_GB50;
wire R5C8_GB10;
wire R16C24_GB50;
wire R26C38_GB20;
wire R10C31_C6;
wire R28C31_Q0;
wire R14C36_GB10;
wire R8C37_GT10;
wire R4C34_GBO0;
wire R5C25_GB50;
wire R11C32_GB20;
wire R28C31_W13;
wire R22C29_GB50;
wire R2C28_GB50;
wire R23C13_GB60;
wire R11C7_GBO0;
wire R28C31_E26;
wire R9C14_GB70;
wire R16C43_GBO1;
wire R28C22_E81;
wire R28C28_S10;
wire R6C14_GB00;
wire R11C14_GT00;
wire R10C34_W21;
wire R15C4_GBO1;
wire R26C36_GB10;
wire R27C35_GB30;
wire R28C31_N21;
wire R6C33_GT10;
wire R4C1_GT00;
wire R5C23_GT00;
wire R28C19_S12;
wire R3C4_GB70;
wire R12C17_GB00;
wire R20C24_GB00;
wire R15C18_GB50;
wire R28C22_N83;
wire R28C13_Q6;
wire R27C6_GB70;
wire R10C7_S22;
wire R28C25_W23;
wire R28C34_CLK2;
wire R6C37_GB10;
wire R7C4_GB40;
wire R27C40_GB40;
wire R1C47_F2;
wire R10C10_E21;
wire R2C40_GB50;
wire R7C15_GB70;
wire R10C13_X07;
wire R27C2_GT10;
wire R21C36_GB30;
wire R28C10_X04;
wire R13C42_GB60;
wire R28C40_D6;
wire R2C25_GB30;
wire R9C18_GBO1;
wire R8C42_GT00;
wire R10C37_EW10;
wire R22C9_GB10;
wire R7C35_GB20;
wire R16C39_GB10;
wire R16C12_GT00;
wire R7C29_GB00;
wire R6C10_GB00;
wire R4C20_GB60;
wire R17C14_GB50;
wire R28C28_CLK2;
wire R15C20_GT10;
wire R28C13_B1;
wire R27C13_GB30;
wire R23C6_GB10;
wire R12C32_GT10;
wire R8C46_GBO0;
wire R20C13_GB00;
wire R10C40_A4;
wire R1C47_C5;
wire R16C3_GBO0;
wire R6C43_GB10;
wire R1C32_W83;
wire R6C28_GB20;
wire R20C21_GB60;
wire R2C4_GBO1;
wire R23C14_GB10;
wire R7C37_GB70;
wire R28C25_D5;
wire R1C47_C2;
wire R28C7_N82;
wire R28C13_Q3;
wire R10C13_Q5;
wire R23C13_GB00;
wire R2C42_GB50;
wire R10C16_W80;
wire R8C20_GB10;
wire R6C37_GB60;
wire R15C15_GBO0;
wire R21C13_GB20;
wire R26C13_GB30;
wire R27C36_GB10;
wire R24C32_GB20;
wire R9C20_GBO1;
wire R3C22_GB70;
wire R17C14_GB00;
wire R10C10_S83;
wire R28C46_CLK1;
wire R22C30_GB00;
wire R8C32_GB00;
wire R16C40_GB00;
wire R15C23_GBO1;
wire R1C28_SEL3;
wire R9C29_GB70;
wire R21C3_GB70;
wire R22C26_GB50;
wire R5C34_GT10;
wire R16C39_GB00;
wire R21C46_GB40;
wire R1C32_D7;
wire R28C7_N24;
wire R14C34_GB00;
wire R17C4_GT00;
wire R10C16_E80;
wire R10C27_E25;
wire R10C22_W80;
wire R27C33_GT10;
wire R20C25_SPINE19;
wire R15C21_GB70;
wire R18C18_GB70;
wire R18C23_GB70;
wire R14C9_GB60;
wire R29C28_X03;
wire R2C13_GB00;
wire R18C44_GB30;
wire R10C30_D6;
wire R2C23_GBO0;
wire R16C13_GBO1;
wire R22C43_GB30;
wire R6C15_GT10;
wire R14C2_GB10;
wire R10C7_N80;
wire R23C39_GT00;
wire R7C23_GBO1;
wire R16C38_GT10;
wire R25C45_GT00;
wire R26C5_GB70;
wire R24C34_GBO0;
wire R28C46_F1;
wire R7C12_GB40;
wire R4C6_GBO1;
wire R14C33_GB70;
wire R22C32_GB70;
wire R12C43_GT10;
wire R24C14_GB10;
wire R28C37_A7;
wire R1C32_A2;
wire R23C2_GB40;
wire R21C35_GB50;
wire R27C29_GT00;
wire R3C34_GBO0;
wire R8C32_GB60;
wire R22C18_GB60;
wire R5C18_GB20;
wire R28C22_N20;
wire R10C29_CLK0;
wire R10C40_C1;
wire R6C19_GB60;
wire R25C44_GT10;
wire R4C39_GB10;
wire R21C31_GB70;
wire R15C1_GT00;
wire R14C44_GB00;
wire R17C24_GB30;
wire R9C25_GBO0;
wire R15C46_GB20;
wire R28C46_A7;
wire R2C23_GT00;
wire R9C7_GB20;
wire R7C14_GB60;
wire R28C19_F7;
wire R28C31_A7;
wire R21C38_GB10;
wire R23C6_GB60;
wire R18C2_GB10;
wire R14C42_GBO1;
wire R20C34_GT10;
wire R16C3_GB40;
wire R28C46_Q6;
wire R14C24_GT00;
wire R23C23_GT10;
wire R4C9_GB50;
wire R11C5_GBO1;
wire R2C10_GB20;
wire R26C35_GB00;
wire R12C31_GB00;
wire R28C28_S27;
wire R10C27_A4;
wire R12C43_GB30;
wire R24C42_GB60;
wire R28C16_C1;
wire R29C28_Q5;
wire R24C40_GT00;
wire R8C38_GB30;
wire R7C22_GB70;
wire R9C12_GB70;
wire R17C13_GB30;
wire R4C15_GB20;
wire R12C24_GB30;
wire R13C39_GB20;
wire R15C5_GB00;
wire R13C41_GB40;
wire R10C22_C3;
wire R28C7_W13;
wire R12C11_GB10;
wire R12C10_GBO1;
wire R28C40_B3;
wire R12C13_GB10;
wire R2C25_GB20;
wire R10C10_E20;
wire R7C16_GB50;
wire R14C6_GB60;
wire R10C28_B4;
wire R14C45_GB60;
wire R28C22_W80;
wire R7C14_GBO1;
wire R16C33_GT00;
wire R6C17_GB60;
wire R8C43_GB50;
wire R7C36_GB60;
wire R27C35_GB60;
wire R28C43_W26;
wire R27C19_GB60;
wire R12C39_GB00;
wire R23C32_GT00;
wire R24C42_GB30;
wire R9C25_GBO1;
wire R28C34_D5;
wire R2C5_GB40;
wire R22C39_GB00;
wire R12C4_GB40;
wire R10C25_X07;
wire R3C29_GB20;
wire R14C35_GBO1;
wire R1C47_S83;
wire R21C5_GB60;
wire R24C4_GBO1;
wire R6C15_GBO0;
wire R11C38_GB10;
wire R14C46_GB50;
wire R18C24_GB10;
wire R28C10_Q4;
wire R5C26_GB20;
wire R20C9_GB40;
wire R28C13_SEL5;
wire R10C43_Q5;
wire R26C34_GB10;
wire R22C18_GB70;
wire R27C11_GB70;
wire R2C44_GB30;
wire R8C17_GT10;
wire R20C31_GBO1;
wire R18C43_GT00;
wire R28C40_W23;
wire R7C45_GB60;
wire R2C44_SPINE0;
wire R24C11_GB20;
wire R14C41_GT00;
wire R20C28_GB60;
wire R1C32_X08;
wire R22C45_GB30;
wire R5C38_GB30;
wire R28C25_A0;
wire R29C28_W26;
wire R20C9_GB70;
wire R12C41_GBO0;
wire R13C38_GB40;
wire R18C27_GT10;
wire R2C39_GB10;
wire R28C16_Q1;
wire R5C17_GB00;
wire R3C27_GB60;
wire R20C41_GT00;
wire R22C4_GT00;
wire R15C13_GB50;
wire R11C1_GBO0;
wire R8C29_GB30;
wire R16C43_GBO0;
wire R14C43_GB60;
wire R1C1_E23;
wire R28C16_N27;
wire R10C27_CLK1;
wire R9C26_GB30;
wire R2C46_GB10;
wire R10C34_N24;
wire R28C16_CLK0;
wire R10C10_SEL4;
wire R28C28_W27;
wire R16C44_GB50;
wire R10C40_S83;
wire R11C43_GB20;
wire R5C32_GB70;
wire R28C13_E13;
wire R17C32_GB70;
wire R21C9_GT00;
wire R11C22_GB50;
wire R22C7_GT00;
wire R10C26_N21;
wire R12C1_GT00;
wire R12C8_GT00;
wire R4C18_GB40;
wire R7C33_GT00;
wire R15C20_GBO1;
wire R3C45_GBO1;
wire R28C10_S12;
wire R28C22_E82;
wire R13C5_GB70;
wire R11C28_GB20;
wire R12C17_GB40;
wire R4C36_GB00;
wire R14C39_GB20;
wire R22C32_GB30;
wire R25C33_GB60;
wire R12C7_GB60;
wire R9C35_GT10;
wire R16C45_GB00;
wire R1C47_B2;
wire R18C30_GBO0;
wire R10C37_E11;
wire R2C11_GB70;
wire R3C30_GB60;
wire R27C38_GBO1;
wire R18C33_GB70;
wire R10C25_W81;
wire R10C40_S27;
wire R14C12_GB40;
wire R7C23_GT00;
wire R28C43_S23;
wire R12C30_GB00;
wire R10C28_W21;
wire R6C11_GB30;
wire R10C25_S24;
wire R5C23_GBO0;
wire R10C28_W25;
wire R22C17_GBO1;
wire R25C27_GB20;
wire R26C34_GB40;
wire R15C35_GB50;
wire R10C13_D4;
wire R2C20_GB60;
wire R2C7_SPINE13;
wire R11C13_GB00;
wire R15C7_GB20;
wire R18C20_GBO1;
wire R27C15_GB50;
wire R4C23_GB00;
wire R15C12_GB70;
wire R3C36_GBO0;
wire R7C32_GB40;
wire R28C10_W82;
wire R22C15_GT00;
wire R13C17_GB00;
wire R2C7_GB20;
wire R5C15_GT00;
wire R8C31_GT10;
wire R15C36_GT10;
wire R22C22_GB30;
wire R22C20_GB50;
wire R8C35_GB00;
wire R13C35_GB00;
wire R24C39_GB20;
wire R15C43_GB60;
wire R23C41_GB70;
wire R10C27_N11;
wire R28C10_S20;
wire R10C30_W12;
wire R3C12_GB10;
wire R18C22_GB20;
wire R5C26_GB60;
wire R28C13_C5;
wire R28C10_CLK2;
wire R1C1_F7;
wire R10C25_D6;
wire R16C24_GT10;
wire R4C36_GB30;
wire R10C30_F4;
wire R28C22_C0;
wire R28C25_F2;
wire R9C7_GB40;
wire R28C19_S81;
wire R22C37_GB60;
wire R28C22_W13;
wire R23C20_GB50;
wire R10C37_S82;
wire R13C38_GT10;
wire R8C11_GB70;
wire R12C22_GB00;
wire R15C39_GBO0;
wire R5C45_GBO0;
wire R4C3_GB70;
wire R10C22_W12;
wire R28C25_E24;
wire R24C28_GB70;
wire R3C35_GB60;
wire R28C46_Q4;
wire R10C31_W24;
wire R28C43_W10;
wire R3C19_GT10;
wire R17C45_GB50;
wire R29C28_S27;
wire R7C42_GB10;
wire R8C27_GT10;
wire R4C25_GB20;
wire R10C29_E25;
wire R18C36_GB30;
wire R20C39_GT00;
wire R10C7_N24;
wire R2C4_GB60;
wire R15C10_GB20;
wire R10C40_D0;
wire R17C40_GB10;
wire R26C28_GB50;
wire R10C28_Q4;
wire R16C41_GT10;
wire R27C16_GB10;
wire R10C16_F6;
wire R28C4_SN10;
wire R10C40_S81;
wire R21C41_GB40;
wire R16C36_GB40;
wire R17C37_GB60;
wire R27C22_GT00;
wire R15C27_GT00;
wire R18C43_GBO0;
wire R10C28_EW20;
wire R28C28_E24;
wire R17C16_GT00;
wire R13C40_GT00;
wire R28C37_X05;
wire R1C1_N26;
wire R10C29_E22;
wire R26C20_GB60;
wire R10C25_F0;
wire R25C30_GT00;
wire R28C37_N20;
wire R1C47_E25;
wire R18C10_GBO1;
wire R11C16_GT10;
wire R11C21_GB70;
wire R25C20_GB00;
wire R28C34_EW10;
wire R20C12_GT00;
wire R6C19_GT10;
wire R16C44_GT10;
wire R15C24_GB00;
wire R12C45_GBO1;
wire R10C29_SPINE28;
wire R18C28_GT00;
wire R15C34_GT00;
wire R14C19_GBO1;
wire R10C29_X08;
wire R4C37_GB60;
wire R27C9_GB30;
wire R5C16_GT00;
wire R2C44_GBO1;
wire R1C28_W22;
wire R24C42_GT00;
wire R9C45_GB10;
wire R26C37_GB60;
wire R2C9_GB10;
wire R7C20_GB40;
wire R21C13_GB60;
wire R26C30_GB10;
wire R20C43_SPINE25;
wire R21C16_GB60;
wire R11C2_GBO0;
wire R24C37_GB40;
wire R4C11_GB30;
wire R11C39_GBO0;
wire R2C7_GB40;
wire R10C30_Q4;
wire R25C19_GB20;
wire R24C6_GB20;
wire R23C22_GT00;
wire R10C30_C6;
wire R11C23_GB60;
wire R20C44_GT00;
wire R4C16_GB10;
wire R13C43_GBO0;
wire R25C22_GB40;
wire R18C36_GB40;
wire R23C40_GB50;
wire R12C46_GT00;
wire R13C13_GB10;
wire R23C5_GBO1;
wire R15C41_GB70;
wire R14C39_GB00;
wire R10C29_E81;
wire R28C16_CLK2;
wire R8C22_GB20;
wire R7C5_GB60;
wire R26C25_GBO1;
wire R20C24_GB40;
wire R10C28_X04;
wire R15C41_GB20;
wire R28C34_N22;
wire R10C16_F5;
wire R25C46_GB60;
wire R14C31_GB10;
wire R28C22_N12;
wire R28C19_C6;
wire R17C40_GB40;
wire R21C27_GB10;
wire R15C21_GB60;
wire R27C43_GB00;
wire R9C36_GT10;
wire R22C11_GB60;
wire R1C28_LSR1;
wire R10C28_UNK121;
wire R10C29_W80;
wire R10C40_X06;
wire R28C4_C7;
wire R24C26_GT10;
wire R24C31_GB30;
wire R10C7_W83;
wire R25C43_GB50;
wire R15C38_GB40;
wire R6C34_GB20;
wire R22C30_GB10;
wire R10C30_N82;
wire R22C21_GB20;
wire R21C29_GBO1;
wire R21C40_GB60;
wire R17C3_GT00;
wire R18C45_GBO0;
wire R28C31_A1;
wire R21C26_GB10;
wire R18C41_GB40;
wire R28C46_S26;
wire R10C13_C2;
wire R28C37_N13;
wire R12C7_GB20;
wire R12C36_GT10;
wire R24C36_GT10;
wire R28C34_S24;
wire R29C28_B1;
wire R3C30_GB00;
wire R2C40_GB20;
wire R14C20_GBO0;
wire R21C38_GBO1;
wire R24C7_GT10;
wire R3C32_GB40;
wire R6C15_GB70;
wire R17C31_GB30;
wire R16C14_GB40;
wire R7C34_GB20;
wire R16C41_GB50;
wire R10C29_N11;
wire R10C25_S81;
wire R28C22_D3;
wire R8C18_GBO1;
wire R13C15_GB50;
wire R3C13_GB00;
wire R16C7_GB00;
wire R6C29_GB50;
wire R4C39_GB30;
wire R12C29_GT10;
wire R10C37_CE2;
wire R8C39_GB30;
wire R11C17_GT00;
wire R10C43_S25;
wire R1C28_N26;
wire R10C10_S82;
wire R6C17_GB70;
wire R2C43_GB60;
wire R14C25_GB70;
wire R8C40_GB50;
wire R15C42_GB50;
wire R1C32_W24;
wire R7C7_GB00;
wire R20C18_GB00;
wire R12C13_GBO0;
wire R18C35_GBO1;
wire R14C12_GB60;
wire R3C40_GT00;
wire R7C28_GB30;
wire R18C37_GBO1;
wire R10C19_E27;
wire R28C7_A3;
wire R14C4_GT10;
wire R22C45_GB50;
wire R17C1_GBO0;
wire R18C3_GB60;
wire R28C16_W10;
wire R10C29_SPINE27;
wire R23C35_GT00;
wire R15C7_GBO0;
wire R13C45_GB50;
wire R24C33_GB30;
wire R2C37_SPINE3;
wire R14C36_GB50;
wire R20C35_SPINE25;
wire R26C46_GB40;
wire R28C19_CE2;
wire R14C13_GB00;
wire R20C9_GT10;
wire R26C10_GB20;
wire R1C1_N27;
wire R10C31_W21;
wire R28C46_N20;
wire R28C34_C5;
wire R16C21_GB70;
wire R11C32_GB00;
wire R13C12_GT10;
wire R12C29_GB00;
wire R6C40_GB50;
wire R23C3_GBO0;
wire R2C30_GBO0;
wire R6C12_GT00;
wire R15C24_GT10;
wire R4C38_GB60;
wire R13C29_GB10;
wire R16C38_GB60;
wire R12C28_GB00;
wire R10C31_S23;
wire R28C7_N83;
wire R3C31_GB50;
wire R23C27_GB20;
wire R28C40_F4;
wire R13C17_GT10;
wire R3C36_GB10;
wire R10C28_UNK128;
wire R5C36_GBO1;
wire R9C17_GB40;
wire R6C35_GB10;
wire R28C4_Q3;
wire R14C27_GB70;
wire R6C46_GBO1;
wire R14C20_GB20;
wire R21C3_GB30;
wire R27C4_GB10;
wire R21C40_GB20;
wire R10C28_W10;
wire R28C13_E26;
wire R6C41_GT10;
wire R3C20_GB60;
wire R11C13_GB70;
wire R26C26_GB60;
wire R28C4_SEL2;
wire R28C22_X03;
wire R21C14_GBO0;
wire R28C37_D2;
wire R20C35_GB70;
wire R1C28_F2;
wire R16C4_GBO0;
wire R8C20_GB40;
wire R10C13_F1;
wire R2C30_GT10;
wire R27C21_GBO0;
wire R1C28_B0;
wire R28C13_S82;
wire R26C11_GB20;
wire R14C35_GB00;
wire R17C43_GB70;
wire R28C37_E12;
wire R17C34_GT10;
wire R28C43_F3;
wire R24C1_GBO0;
wire R1C28_E20;
wire R12C10_GBO0;
wire R16C24_GBO0;
wire R11C13_GBO0;
wire R10C10_CLK0;
wire R28C10_LSR2;
wire R5C35_GB40;
wire R5C8_GT10;
wire R20C42_GBO1;
wire R10C30_EW20;
wire R27C17_GB10;
wire R14C12_GT00;
wire R27C38_GT10;
wire R3C45_GB40;
wire R20C28_GB50;
wire R20C32_GB70;
wire R2C23_GB20;
wire R14C10_GB20;
wire R10C7_W20;
wire R3C6_GB40;
wire R18C26_GB30;
wire R14C10_GT10;
wire R13C43_GT00;
wire R26C32_GB00;
wire R10C25_E27;
wire R10C34_N83;
wire R15C44_GT10;
wire R28C16_S22;
wire R27C9_GB70;
wire R2C36_GB50;
wire R28C25_B0;
wire R28C25_E82;
wire R20C35_GT00;
wire R20C43_GT00;
wire R9C15_GB50;
wire R3C32_GB50;
wire R1C32_D3;
wire R21C1_GT00;
wire R10C29_W23;
wire R18C12_GB10;
wire R7C46_GB30;
wire R2C37_GB70;
wire R4C15_GB00;
wire R9C9_GB10;
wire R4C9_GBO0;
wire R28C43_N12;
wire R18C46_GB70;
wire R5C26_GBO1;
wire R8C15_GB60;
wire R25C6_GBO0;
wire R12C38_GB40;
wire R11C34_GB30;
wire R28C46_X04;
wire R16C24_GB60;
wire R10C29_A3;
wire R25C5_GB20;
wire R15C40_GB50;
wire R12C16_GB70;
wire R20C14_GT00;
wire R26C23_GB50;
wire R10C34_B3;
wire R28C22_C5;
wire R4C7_GBO1;
wire R27C23_GB50;
wire R28C10_W27;
wire R17C38_GB40;
wire R4C9_GBO1;
wire R26C28_GB70;
wire R6C6_GB40;
wire R10C19_E25;
wire R12C32_GBO0;
wire R28C22_B1;
wire R22C21_GT00;
wire R24C15_GB60;
wire R16C11_GT00;
wire R5C39_GBO0;
wire R2C38_GB40;
wire R1C32_E24;
wire R25C16_GB60;
wire R10C37_S11;
wire R10C22_Q1;
wire R20C23_GB00;
wire R2C41_GB10;
wire R8C18_GB40;
wire R15C44_GB70;
wire R27C27_GT00;
wire R16C32_GBO0;
wire R16C12_GBO1;
wire R13C36_GBO0;
wire R24C10_GB00;
wire R24C29_GB00;
wire R4C40_GB00;
wire R14C10_GB10;
wire R25C38_GB10;
wire R17C35_GB00;
wire R5C9_GT00;
wire R28C10_F5;
wire R24C20_GBO0;
wire R6C21_GBO1;
wire R6C16_GBO0;
wire R10C26_C1;
wire R10C27_E11;
wire R10C29_F2;
wire R11C15_GBO1;
wire R15C18_GBO1;
wire R14C3_GB20;
wire R13C33_GB70;
wire R24C16_GT10;
wire R23C4_GB10;
wire R20C31_GT10;
wire R24C16_GB60;
wire R11C46_GB20;
wire R10C40_N11;
wire R9C12_GT10;
wire R23C40_GBO0;
wire R20C3_GB60;
wire R10C28_N83;
wire R23C21_GB30;
wire R22C5_GB60;
wire R8C21_GB20;
wire R10C31_N21;
wire R27C5_GB60;
wire R9C2_GBO0;
wire R27C14_GB50;
wire R11C6_GT10;
wire R3C46_GB30;
wire R3C6_GT00;
wire R5C21_GB20;
wire R2C42_GBO0;
wire R22C35_GB50;
wire R10C27_E12;
wire R8C13_GB50;
wire R11C46_GT00;
wire R11C9_GB00;
wire R16C4_GB60;
wire R25C26_GB00;
wire R12C26_GB70;
wire R27C22_GB60;
wire R14C39_GB10;
wire R26C40_GT00;
wire R28C4_S24;
wire R2C20_GB40;
wire R22C22_GB70;
wire R23C15_GB10;
wire R20C19_GB20;
wire R10C10_B5;
wire R13C24_GT00;
wire R9C12_GB30;
wire R16C19_GB00;
wire R3C37_GB00;
wire R12C7_GB50;
wire R10C27_UNK126;
wire R22C23_GB00;
wire R16C17_GBO0;
wire R28C31_F3;
wire R5C40_GT00;
wire R16C26_GB20;
wire R6C33_GB50;
wire R18C21_GT00;
wire R25C39_GBO0;
wire R24C25_GB00;
wire R28C10_N11;
wire R11C30_GT10;
wire R29C28_F6;
wire R17C35_GT10;
wire R2C46_GB00;
wire R10C19_S12;
wire R4C5_GB00;
wire R8C9_GB20;
wire R10C13_D3;
wire R10C28_C2;
wire R1C28_S82;
wire R11C17_GB50;
wire R10C40_A6;
wire R25C15_GB00;
wire R8C16_GBO0;
wire R23C27_GB00;
wire R28C13_A3;
wire R4C40_GB10;
wire R24C3_GB00;
wire R28C43_N24;
wire R20C16_GB40;
wire R28C40_Q0;
wire R7C15_GB20;
wire R13C24_GB60;
wire R22C43_GB10;
wire R13C2_GB00;
wire R3C38_GT10;
wire R10C22_F3;
wire R1C29_F6;
wire R26C31_GB30;
wire R24C22_GB20;
wire R10C34_D2;
wire R26C46_GB60;
wire R10C28_SPINE21;
wire R23C11_GT00;
wire R12C46_GBO0;
wire R23C35_GB50;
wire R20C31_GB70;
wire R8C4_GB40;
wire R10C34_Q4;
wire R4C13_GB00;
wire R16C21_GB20;
wire R5C39_GB40;
wire R7C37_GBO1;
wire R18C28_GB00;
wire R17C36_GBO1;
wire R27C32_GB70;
wire R28C31_LSR2;
wire R28C10_E11;
wire R15C22_GB60;
wire R10C16_Q1;
wire R17C33_GB60;
wire R16C1_GBO0;
wire R28C13_N27;
wire R8C43_GB20;
wire R27C10_GB60;
wire R16C32_GB30;
wire R28C25_N24;
wire R2C21_GBO1;
wire R4C4_GB60;
wire R10C28_N27;
wire R9C43_GT00;
wire R25C31_GB70;
wire R5C26_GBO0;
wire R12C20_GB00;
wire R14C2_GT10;
wire R20C28_GB30;
wire R9C45_GB20;
wire R20C18_GB40;
wire R8C44_GB70;
wire R5C26_GB10;
wire R5C38_GT00;
wire R2C9_GB70;
wire R21C11_GB40;
wire R4C44_GB50;
wire R25C33_GB30;
wire R4C36_GBO1;
wire R10C30_S22;
wire R22C11_GB10;
wire R10C22_LSR2;
wire R20C37_GB00;
wire R10C30_CLK1;
wire R28C10_N80;
wire R14C36_GB20;
wire R11C28_GT00;
wire R5C43_GBO1;
wire R17C28_GB00;
wire R28C22_A1;
wire R16C39_GBO1;
wire R25C31_GB00;
wire R11C10_GT00;
wire R20C19_GT10;
wire R12C6_GBO0;
wire R1C47_E26;
wire R14C43_GBO1;
wire R2C15_GT00;
wire R9C10_GB10;
wire R10C26_N20;
wire R11C17_GB20;
wire R15C36_GB30;
wire R13C20_GB60;
wire R27C22_GT10;
wire R14C41_GB40;
wire R18C41_GB00;
wire R15C32_GB20;
wire R28C7_E23;
wire R25C5_GT10;
wire R28C22_F2;
wire R10C30_UNK121;
wire R23C40_GB40;
wire R13C24_GB70;
wire R3C41_GT10;
wire R24C2_GT10;
wire R17C35_GB70;
wire R3C3_GB30;
wire R10C27_Q1;
wire R4C21_GT10;
wire R3C40_GT10;
wire R26C7_GB30;
wire R18C20_GB30;
wire R29C28_S13;
wire R5C14_GB50;
wire R8C32_GB70;
wire R28C25_X06;
wire R14C27_GT00;
wire R10C29_C2;
wire R23C5_GB60;
wire R28C4_S13;
wire R10C22_E81;
wire R5C46_GB60;
wire R22C40_GB20;
wire R1C47_S22;
wire R2C3_GB10;
wire R1C1_W26;
wire R24C44_GB50;
wire R1C47_N23;
wire R11C7_GB30;
wire R15C16_GB70;
wire R15C31_GB70;
wire R10C26_B3;
wire R10C29_X05;
wire R8C20_GB60;
wire R24C18_GB40;
wire R9C22_GT00;
wire R3C14_GBO1;
wire R24C28_GB50;
wire R15C37_GB70;
wire R28C46_N13;
wire R23C16_GB20;
wire R10C13_X05;
wire R28C40_W12;
wire R16C36_GB20;
wire R15C27_GB30;
wire R28C37_D3;
wire R6C8_GBO1;
wire R9C6_GB50;
wire R29C28_W21;
wire R18C6_GB20;
wire R2C38_GB10;
wire R3C46_GBO0;
wire R11C35_GB60;
wire R7C31_GB50;
wire R2C30_GB10;
wire R22C45_GT10;
wire R7C26_GB50;
wire R5C32_GBO0;
wire R10C10_N11;
wire R28C19_D1;
wire R15C23_GB40;
wire R22C6_GBO1;
wire R11C6_GB10;
wire R20C19_GB30;
wire R4C29_GBO0;
wire R9C12_GB60;
wire R28C43_SEL3;
wire R12C25_GB30;
wire R21C12_GB50;
wire R28C46_E13;
wire R3C37_GB40;
wire R22C29_GB60;
wire R14C14_GT10;
wire R10C30_SPINE2;
wire R23C31_GT00;
wire R5C12_GB70;
wire R5C33_GB70;
wire R24C31_GB40;
wire R17C33_GBO1;
wire R28C19_B1;
wire R18C13_GB10;
wire R22C43_GB00;
wire R29C28_N83;
wire R26C4_GB10;
wire R25C20_GB30;
wire R9C41_GB40;
wire R10C29_N13;
wire R4C29_GB20;
wire R12C26_GT00;
wire R25C20_GB20;
wire R13C30_GT10;
wire R17C11_GB60;
wire R1C47_W24;
wire R10C22_C0;
wire R18C14_GB00;
wire R1C28_X07;
wire R28C43_W24;
wire R28C31_CE1;
wire R28C37_F0;
wire R26C24_GT00;
wire R6C33_GBO0;
wire R2C35_SPINE5;
wire R21C10_GB30;
wire R3C44_GT10;
wire R25C12_GB10;
wire R4C45_GBO0;
wire R6C24_GB30;
wire R5C34_GB60;
wire R27C24_GB50;
wire R10C43_S83;
wire R11C18_GB10;
wire R25C9_GBO0;
wire R28C40_N83;
wire R5C41_GBO0;
wire R18C33_GB10;
wire R28C40_S22;
wire R5C43_GB70;
wire R23C23_GBO1;
wire R6C9_GB30;
wire R25C18_GB50;
wire R26C12_GB30;
wire R27C37_GB70;
wire R1C1_Q1;
wire R25C33_GB10;
wire R20C26_GB70;
wire R1C47_C0;
wire R10C26_N83;
wire R26C46_GB50;
wire R25C29_GBO1;
wire R25C29_GT00;
wire R28C10_W81;
wire R2C17_GB00;
wire R28C22_N82;
wire R28C34_W26;
wire R10C37_CLK2;
wire R25C45_GB40;
wire R13C10_GB20;
wire R11C5_GT00;
wire R16C21_GB40;
wire R9C9_GB40;
wire R11C3_GB10;
wire R25C18_GB70;
wire R4C32_GB20;
wire R8C33_GT10;
wire R11C13_GB10;
wire R24C4_GT00;
wire R17C17_GB00;
wire R26C24_GBO0;
wire R27C14_GB20;
wire R20C34_GB10;
wire R7C10_GB00;
wire R9C25_GB30;
wire R8C13_GBO1;
wire R7C9_GT10;
wire R2C28_GB30;
wire R6C12_GBO0;
wire R10C40_CE1;
wire R12C12_GBO1;
wire R17C32_GBO1;
wire R28C46_A3;
wire R2C3_GB40;
wire R14C31_GT00;
wire R11C12_GB40;
wire R9C28_GB70;
wire R23C25_GT00;
wire R10C31_A5;
wire R7C17_GT10;
wire R10C27_SEL5;
wire R4C39_GBO1;
wire R12C34_GB00;
wire R9C5_GT10;
wire R13C9_GB50;
wire R7C39_GB20;
wire R28C10_S24;
wire R28C25_A7;
wire R4C3_GT00;
wire R25C23_GB10;
wire R23C34_GB60;
wire R28C16_W25;
wire R4C46_GB20;
wire R6C19_GBO1;
wire R3C44_GB20;
wire R17C29_GB50;
wire R28C46_W10;
wire R22C32_GB60;
wire R10C31_LSR1;
wire R28C13_E24;
wire R13C37_GB20;
wire R10C43_X05;
wire R10C40_X04;
wire R28C19_Q0;
wire R28C16_CE0;
wire R3C8_GB60;
wire R15C2_GB00;
wire R20C33_GB30;
wire R10C19_D7;
wire R10C22_N26;
wire R23C16_GB50;
wire R14C3_GB70;
wire R17C1_GT10;
wire R10C28_E82;
wire R4C10_GB20;
wire R10C29_N81;
wire R27C18_GB60;
wire R5C38_GB60;
wire R28C28_E83;
wire R15C19_GB70;
wire R13C25_GBO1;
wire R20C42_GB70;
wire R15C28_GB40;
wire R23C24_GBO1;
wire R10C27_X03;
wire R2C46_GBO0;
wire R16C5_GT10;
wire R10C29_W20;
wire R1C32_N83;
wire R2C26_GT00;
wire R28C46_W11;
wire R28C46_F0;
wire R8C4_GT00;
wire R25C25_GBO1;
wire R8C29_GT10;
wire R5C16_GB10;
wire R27C23_GB30;
wire R13C27_GB40;
wire R9C36_GB00;
wire R28C31_W24;
wire R18C42_GB50;
wire R12C35_GBO0;
wire R11C33_GB60;
wire R24C44_GBO1;
wire R12C30_GB70;
wire R2C5_GT10;
wire R6C37_GB40;
wire R21C6_GB30;
wire R20C4_GB40;
wire R14C28_GB50;
wire R1C28_F5;
wire R21C32_GT00;
wire R24C37_GB70;
wire R14C14_GBO0;
wire R5C35_GB50;
wire R10C28_S25;
wire R11C8_GB10;
wire R4C32_GB60;
wire R23C35_GBO0;
wire R23C27_GB70;
wire R10C31_X02;
wire R3C39_GBO1;
wire R7C24_GB00;
wire R26C31_GBO0;
wire R10C31_X07;
wire R10C31_C4;
wire R20C16_GB20;
wire R3C23_GB00;
wire R25C18_GB00;
wire R6C33_GB70;
wire R7C16_GBO1;
wire R28C43_D5;
wire R20C38_GB30;
wire R18C43_GB40;
wire R6C22_GBO1;
wire R17C7_GB10;
wire R1C32_E81;
wire R5C37_GB60;
wire R20C6_GB40;
wire R10C7_N13;
wire R13C4_GB50;
wire R21C5_GB20;
wire R12C15_GT00;
wire R10C27_S23;
wire R18C38_GB70;
wire R25C13_GB10;
wire R10C31_A1;
wire R7C17_GB50;
wire R23C28_GB40;
wire R22C3_GB50;
wire R5C15_GB60;
wire R18C23_GB00;
wire R21C26_GBO0;
wire R27C6_GB40;
wire R28C25_N23;
wire R5C35_GT00;
wire R18C27_GB50;
wire R25C37_GB40;
wire R8C9_GB60;
wire R10C26_CLK2;
wire R7C8_GB50;
wire R15C11_GB10;
wire R21C37_GB00;
wire R28C16_X04;
wire R11C20_GB10;
wire R11C36_GB60;
wire R28C37_S80;
wire R15C4_GB60;
wire R20C9_GB00;
wire R2C33_GBO0;
wire R10C27_D6;
wire R28C13_W23;
wire R17C42_GB20;
wire R10C40_C5;
wire R10C27_X08;
wire R10C26_S26;
wire R10C10_W20;
wire R27C7_GB40;
wire R24C31_GBO1;
wire R10C40_W82;
wire R28C7_E11;
wire R26C22_GB20;
wire R28C4_N11;
wire R10C25_E24;
wire R2C26_GB40;
wire R26C26_GB10;
wire R14C16_GB20;
wire R15C15_GB50;
wire R28C13_S23;
wire R22C22_GBO1;
wire R28C4_LSR0;
wire R13C14_GB50;
wire R28C37_B2;
wire R24C43_GT10;
wire R20C22_GB40;
wire R11C10_GB10;
wire R10C16_SEL7;
wire R2C4_GB10;
wire R1C28_Q0;
wire R10C13_W83;
wire R7C4_GT00;
wire R6C1_GBO1;
wire R23C45_GBO0;
wire R20C3_GBO0;
wire R3C29_GBO1;
wire R1C32_F0;
wire R3C8_GBO0;
wire R10C19_X04;
wire R5C6_GB50;
wire R5C4_GB00;
wire R15C43_GB00;
wire R21C39_GB60;
wire R28C10_C5;
wire R10C26_W83;
wire R2C40_GB60;
wire R21C43_GB20;
wire R14C39_GB60;
wire R27C11_GT00;
wire R16C13_GT00;
wire R12C19_GB00;
wire R18C22_GB50;
wire R4C9_GB00;
wire R11C28_GB00;
wire R20C39_GB60;
wire R20C6_GT10;
wire R25C30_GB10;
wire R10C10_S11;
wire R12C28_GT00;
wire R11C45_GT00;
wire R16C3_GT00;
wire R10C30_S20;
wire R21C18_GB30;
wire R15C16_GBO1;
wire R22C2_GB70;
wire R28C46_D5;
wire R17C45_GBO1;
wire R28C10_N82;
wire R6C8_GB10;
wire R26C28_GB40;
wire R25C43_GB30;
wire R11C13_GB30;
wire R9C31_GB40;
wire R11C26_GT00;
wire R10C34_C1;
wire R20C7_GT10;
wire R18C6_GT00;
wire R1C1_W13;
wire R13C32_GT00;
wire R28C10_N24;
wire R10C28_D4;
wire R10C28_SEL0;
wire R2C32_GB50;
wire R9C32_GB00;
wire R17C39_GB00;
wire R26C2_GB50;
wire R24C33_GB60;
wire R5C37_GB20;
wire R18C32_GB20;
wire R2C10_GBO0;
wire R10C40_X08;
wire R10C22_B3;
wire R28C22_S25;
wire R26C45_GB50;
wire R8C5_GB60;
wire R28C7_W12;
wire R7C16_GB30;
wire R28C28_Q4;
wire R13C22_GB70;
wire R26C20_GB10;
wire R1C28_SN10;
wire R28C31_S27;
wire R6C16_GB30;
wire R27C5_GBO1;
wire R28C19_E23;
wire R10C7_X02;
wire R21C34_GB40;
wire R28C25_C1;
wire R9C40_GB10;
wire R4C15_GB40;
wire R28C46_N82;
wire R28C43_SEL7;
wire R15C46_GT10;
wire R2C8_GBO1;
wire R2C31_GB70;
wire R11C14_GB50;
wire R1C32_CE2;
wire R28C13_S12;
wire R24C46_GB10;
wire R1C1_E82;
wire R2C21_GB10;
wire R13C10_GBO0;
wire R15C17_GB40;
wire R26C44_GB10;
wire R3C35_GB10;
wire R27C41_GT00;
wire R24C45_GBO0;
wire R10C40_B2;
wire R18C40_GT10;
wire R28C10_N12;
wire R28C25_W20;
wire R25C3_GB50;
wire R2C41_GB70;
wire R2C6_GB70;
wire R26C36_GT10;
wire R3C17_GB00;
wire R23C29_GT10;
wire R28C22_D0;
wire R17C7_GBO0;
wire R15C42_GBO0;
wire R14C19_GB40;
wire R26C35_GB40;
wire R10C25_C4;
wire R14C3_GB40;
wire R3C34_GB20;
wire R4C29_GT00;
wire R23C23_GB40;
wire R15C31_GBO0;
wire R26C3_GB50;
wire R12C39_GB20;
wire R12C40_GB20;
wire R27C13_GB70;
wire R27C31_GB20;
wire R27C46_GB70;
wire R12C15_GB20;
wire R22C26_GBO0;
wire R7C20_GB20;
wire R11C36_GB10;
wire R5C15_GBO1;
wire R5C18_GB10;
wire R12C8_GB70;
wire R12C34_GT10;
wire R20C8_GB20;
wire R3C7_GBO0;
wire R24C20_GB50;
wire R28C19_D0;
wire R5C15_GB00;
wire R14C10_GBO0;
wire R7C32_GBO0;
wire R5C31_GB50;
wire R4C5_GB60;
wire R12C10_GB50;
wire R5C36_GB20;
wire R28C19_LSR1;
wire R10C43_F2;
wire R28C10_SEL5;
wire R27C26_GBO0;
wire R22C37_GB40;
wire R22C13_GB00;
wire R22C12_GB50;
wire R9C27_GT10;
wire R10C22_LSR0;
wire R12C4_GB20;
wire R10C27_SEL4;
wire R11C46_GB30;
wire R28C22_Q3;
wire R11C46_GT10;
wire R8C10_GB50;
wire R16C35_GT10;
wire R11C30_GBO1;
wire R10C10_CE1;
wire R21C23_GB50;
wire R25C40_GB40;
wire R9C19_GT10;
wire R24C14_GBO0;
wire R24C2_GB30;
wire R20C33_SPINE27;
wire R8C4_GT10;
wire R15C45_GB20;
wire R28C10_W11;
wire R4C27_GB20;
wire R10C43_D3;
wire R10C25_S13;
wire R16C22_GB00;
wire R12C24_GB00;
wire R8C17_GB40;
wire R27C24_GBO0;
wire R11C6_GB00;
wire R27C28_GB10;
wire R18C30_GB10;
wire R26C46_GB20;
wire R17C18_GB60;
wire R10C13_D5;
wire R1C47_W27;
wire R5C41_GT10;
wire R6C9_GT00;
wire R9C34_GB40;
wire R13C39_GB60;
wire R16C44_GB70;
wire R3C25_GB20;
wire R28C19_F0;
wire R15C33_GB10;
wire R21C19_GBO0;
wire R15C21_GB00;
wire R21C3_GB40;
wire R18C27_GB60;
wire R1C28_E82;
wire R14C28_GB10;
wire R27C26_GB30;
wire R8C39_GB70;
wire R28C37_A2;
wire R6C12_GB00;
wire R20C9_GB30;
wire R8C8_GB60;
wire R13C1_GBO0;
wire R25C29_GB70;
wire R10C29_W83;
wire R27C3_GB00;
wire R16C38_GBO0;
wire R28C13_E10;
wire R20C21_GT10;
wire R3C46_GB00;
wire R16C13_GB10;
wire R2C37_GB50;
wire R28C10_CE1;
wire R28C31_C4;
wire R23C19_GB50;
wire R15C22_GB70;
wire R5C46_GT10;
wire R11C22_GB20;
wire R17C14_GB70;
wire R10C27_C5;
wire R28C43_B1;
wire R2C35_GBO0;
wire R10C30_A7;
wire R28C19_D3;
wire R17C25_GB20;
wire R14C18_GT10;
wire R13C21_GBO0;
wire R23C17_GB20;
wire R27C13_GBO0;
wire R13C34_GBO1;
wire R1C1_W20;
wire R24C23_GBO1;
wire R3C2_GB60;
wire R16C3_GB10;
wire R10C30_S82;
wire R10C34_Q3;
wire R20C34_GB00;
wire R12C37_GB70;
wire R24C45_GB00;
wire R28C40_W80;
wire R4C41_GT00;
wire R18C33_GB00;
wire R28C25_W21;
wire R28C16_CE2;
wire R10C22_D6;
wire R28C37_F4;
wire R10C27_SEL1;
wire R13C26_GBO1;
wire R24C9_GB20;
wire R2C42_GB40;
wire R14C46_GBO1;
wire R28C34_E11;
wire R26C16_GB50;
wire R20C8_GT10;
wire R6C7_GB10;
wire R14C46_GB00;
wire R20C30_GB10;
wire R11C10_GB70;
wire R24C11_GB60;
wire R12C14_GBO1;
wire R28C31_S25;
wire R24C10_GT10;
wire R10C27_C2;
wire R9C11_GT10;
wire R10C27_UNK127;
wire R2C11_GB60;
wire R8C19_GB40;
wire R26C19_GB40;
wire R5C16_GBO0;
wire R3C38_GB40;
wire R1C28_C4;
wire R10C37_D7;
wire R28C19_D6;
wire R28C10_F7;
wire R17C2_GB70;
wire R10C10_S80;
wire R24C38_GB70;
wire R10C27_W23;
wire R28C40_S82;
wire R13C35_GB70;
wire R10C25_E25;
wire R24C36_GB00;
wire R21C44_GB20;
wire R7C43_GBO1;
wire R16C13_GB20;
wire R26C20_GB30;
wire R6C12_GB10;
wire R8C34_GB50;
wire R3C29_GBO0;
wire R10C13_C5;
wire R27C5_GBO0;
wire R13C1_GBO1;
wire R4C2_GB60;
wire R3C16_GB10;
wire R15C4_GT10;
wire R10C25_D5;
wire R11C5_GB40;
wire R7C42_GB60;
wire R10C7_B4;
wire R10C40_SEL7;
wire R11C1_GT00;
wire R16C26_GB40;
wire R2C33_GB40;
wire R23C5_GB40;
wire R15C46_GBO0;
wire R24C21_GB60;
wire R5C2_GBO0;
wire R6C2_GB00;
wire R14C21_GB40;
wire R27C8_GB30;
wire R10C7_CE1;
wire R21C29_GB40;
wire R27C33_GB10;
wire R13C16_GBO1;
wire R27C25_GB40;
wire R21C31_GBO0;
wire R28C25_W11;
wire R28C37_W21;
wire R13C24_GB20;
wire R28C25_SEL0;
wire R14C34_GB10;
wire R13C35_GT10;
wire R26C19_GB60;
wire R4C41_GB40;
wire R2C21_GBO0;
wire R4C33_GB00;
wire R14C20_GB50;
wire R27C16_GB60;
wire R6C45_GBO1;
wire R29C28_D3;
wire R28C37_Q7;
wire R7C42_GB00;
wire R6C35_GB50;
wire R29C28_F3;
wire R5C15_GB50;
wire R6C34_GBO0;
wire R16C4_GB50;
wire R28C46_E11;
wire R15C11_GBO0;
wire R10C26_N22;
wire R4C13_GT10;
wire R18C26_GB60;
wire R22C41_GB70;
wire R22C20_GB00;
wire R28C46_S80;
wire R27C31_GT00;
wire R2C40_GB00;
wire R28C40_S81;
wire R7C21_GB10;
wire R22C3_GB10;
wire R25C21_GT00;
wire R21C33_GBO0;
wire R12C35_GB00;
wire R23C26_GT00;
wire R20C30_GB20;
wire R5C12_GT10;
wire R23C12_GT00;
wire R2C42_GB20;
wire R22C35_GBO0;
wire R25C42_GB30;
wire R1C28_S13;
wire R26C7_GT10;
wire R5C46_GB00;
wire R28C10_Q2;
wire R7C25_GB60;
wire R28C13_A0;
wire R2C23_GB50;
wire R1C32_N25;
wire R10C28_S83;
wire R28C31_E80;
wire R28C22_F7;
wire R4C39_GB20;
wire R13C22_GB60;
wire R28C4_D2;
wire R28C28_F1;
wire R9C7_GB50;
wire R26C5_GB30;
wire R25C3_GB40;
wire R10C7_B6;
wire R26C18_GB60;
wire R25C20_GT00;
wire R8C10_GBO1;
wire R18C13_GB20;
wire R29C28_E13;
wire R23C23_GB70;
wire R14C28_GB00;
wire R9C2_GB10;
wire R21C11_GB50;
wire R14C27_GBO1;
wire R14C6_GB40;
wire R2C34_GB50;
wire R18C17_GB00;
wire R2C34_GBO0;
wire R23C31_GB70;
wire R15C34_GB70;
wire R11C44_GB60;
wire R16C35_GB40;
wire R28C31_E83;
wire R28C13_LSR2;
wire R7C11_GT10;
wire R8C17_GB50;
wire R6C20_GB50;
wire R26C10_GBO1;
wire R10C34_LSR1;
wire R28C16_E22;
wire R25C38_GBO0;
wire R3C7_GT00;
wire R8C31_GB70;
wire R9C25_GB40;
wire R28C43_Q5;
wire R18C24_GT00;
wire R8C35_GB30;
wire R24C32_GBO0;
wire R12C31_GB60;
wire R10C29_SEL1;
wire R27C41_GB00;
wire R10C28_SN10;
wire R12C17_GB70;
wire R6C18_GB10;
wire R5C40_GB50;
wire R22C11_GBO0;
wire R8C16_GB50;
wire R10C28_X02;
wire R13C13_GB30;
wire R10C31_Q1;
wire R28C25_B7;
wire R23C18_GBO1;
wire R22C10_GB20;
wire R6C2_GB70;
wire R28C43_X08;
wire R24C11_GT00;
wire R22C21_GB60;
wire R13C46_GBO0;
wire R10C22_S22;
wire R25C28_GB00;
wire R16C34_GB70;
wire R24C39_GT10;
wire R1C32_N12;
wire R16C40_GB20;
wire R10C22_E23;
wire R9C21_GB10;
wire R4C13_GB50;
wire R6C28_GB60;
wire R13C4_GB40;
wire R23C34_GT10;
wire R15C18_GB30;
wire R26C38_GT00;
wire R6C36_GBO0;
wire R10C30_F6;
wire R28C37_S13;
wire R18C33_GB30;
wire R18C44_GB00;
wire R28C37_S10;
wire R25C23_GB70;
wire R16C19_GT00;
wire R26C16_GT00;
wire R17C6_GB40;
wire R28C7_C5;
wire R16C42_GT10;
wire R14C19_GT10;
wire R7C11_GB20;
wire R18C21_GB20;
wire R18C8_GB70;
wire R16C29_GB00;
wire R16C19_GB30;
wire R15C3_GBO0;
wire R14C13_GB50;
wire R4C32_GBO0;
wire R26C20_GBO0;
wire R12C32_GB10;
wire R17C34_GB50;
wire R10C16_E81;
wire R10C43_Q2;
wire R10C25_S83;
wire R28C37_SN20;
wire R22C32_GB40;
wire R22C23_GBO0;
wire R4C23_GB50;
wire R13C15_GT00;
wire R6C2_GB30;
wire R5C37_GB70;
wire R27C5_GT10;
wire R18C27_GT00;
wire R14C43_GB30;
wire R10C30_S21;
wire R10C31_EW10;
wire R10C19_W12;
wire R11C7_GT00;
wire R28C16_E81;
wire R28C22_SEL6;
wire R16C46_GB40;
wire R14C36_GBO1;
wire R28C13_W81;
wire R24C9_GBO1;
wire R4C18_GBO1;
wire R6C40_GB60;
wire R17C20_GBO0;
wire R27C25_GT00;
wire R23C39_GB30;
wire R10C19_S25;
wire R27C22_GB50;
wire R27C30_GT10;
wire R6C36_GBO1;
wire R10C27_Q5;
wire R4C35_GB30;
wire R20C26_GB40;
wire R20C8_GB40;
wire R2C46_GB20;
wire R22C30_GB20;
wire R23C32_GBO1;
wire R10C26_D0;
wire R10C28_E20;
wire R10C40_SN20;
wire R28C16_B1;
wire R10C19_C6;
wire R3C5_GBO0;
wire R1C32_N26;
wire R10C40_N82;
wire R10C40_W26;
wire R21C9_GB50;
wire R2C14_GB00;
wire R13C42_GB20;
wire R18C34_GB50;
wire R3C22_GB00;
wire R9C2_GB20;
wire R14C7_GB30;
wire R17C31_GBO1;
wire R18C7_GBO1;
wire R10C27_W11;
wire R1C32_E25;
wire R23C13_GT10;
wire R13C3_GT10;
wire R21C31_GB20;
wire R1C1_X01;
wire R10C7_CLK1;
wire R10C16_X06;
wire R9C22_GB40;
wire R21C23_GB70;
wire R28C34_C4;
wire R13C42_GT00;
wire R26C30_GB40;
wire R26C45_GB70;
wire R4C21_GB60;
wire R10C26_EW10;
wire R28C16_A4;
wire R1C47_N22;
wire R10C37_N83;
wire R10C7_SN10;
wire R18C42_GBO0;
wire R17C33_GB50;
wire R12C44_GB00;
wire R13C12_GT00;
wire R10C34_S27;
wire R18C15_GB70;
wire R29C28_X08;
wire R28C16_S11;
wire R21C26_GB70;
wire R15C14_GT10;
wire R9C32_GBO1;
wire R28C7_W27;
wire R6C35_GB20;
wire R14C22_GT10;
wire R7C40_GB30;
wire R10C19_Q1;
wire R24C43_GBO1;
wire R26C18_GT00;
wire R24C34_GB60;
wire R18C45_GB30;
wire R1C47_X01;
wire R16C2_GB20;
wire R13C44_GBO1;
wire R23C19_GT00;
wire R13C43_GB30;
wire R10C34_E27;
wire R12C4_GB10;
wire R28C13_W10;
wire R25C7_GB40;
wire R4C26_GB10;
wire R8C22_GB50;
wire R17C4_GB30;
wire R14C41_GB60;
wire R10C29_E27;
wire R12C45_GB10;
wire R23C4_GB00;
wire R17C41_GB70;
wire R28C7_B5;
wire R2C17_GBO0;
wire R2C11_GB30;
wire R3C4_GB20;
wire R10C7_C7;
wire R10C22_S26;
wire R27C21_GB00;
wire R18C26_GBO1;
wire R20C22_GB10;
wire R21C12_GB30;
wire R9C11_GB10;
wire R23C43_GB40;
wire R10C43_E25;
wire R18C35_GT00;
wire R27C43_GT00;
wire R8C45_GB30;
wire R10C40_CLK2;
wire R2C35_GB40;
wire R22C33_GT10;
wire R26C8_GB00;
wire R22C29_GB00;
wire R8C33_GB50;
wire R10C26_W24;
wire R16C26_GB30;
wire R16C16_GB20;
wire R10C37_X07;
wire R28C37_W20;
wire R28C28_A1;
wire R28C7_C2;
wire R12C5_GB20;
wire R3C24_GB10;
wire R10C29_W81;
wire R29C28_C2;
wire R7C19_GB00;
wire R9C43_GB20;
wire R1C47_S12;
wire R28C22_E21;
wire R10C22_CE1;
wire R26C29_GT10;
wire R15C2_GB40;
wire R25C6_GB40;
wire R4C34_GB00;
wire R4C36_GB40;
wire R20C41_GB30;
wire R10C31_Q3;
wire R10C30_CE0;
wire R27C11_GBO1;
wire R10C19_S13;
wire R1C1_W22;
wire R28C43_CE0;
wire R4C25_GB50;
wire R10C19_W11;
wire R10C26_F4;
wire R1C32_C1;
wire R14C12_GT10;
wire R27C37_GT10;
wire R22C45_GBO0;
wire R26C15_GB40;
wire R1C1_F2;
wire R24C12_GB10;
wire R10C27_N22;
wire R26C13_GB00;
wire R10C40_LSR2;
wire R16C7_GB40;
wire R28C22_B6;
wire R25C17_GBO1;
wire R26C37_GB00;
wire R13C29_GB40;
wire R28C28_A5;
wire R10C19_A1;
wire R28C34_S23;
wire R9C14_GB00;
wire R23C4_GBO0;
wire R16C45_GBO0;
wire R6C9_GB60;
wire R20C45_GT00;
wire R27C27_GB00;
wire R6C13_GB60;
wire R27C30_GBO1;
wire R28C10_N26;
wire R5C23_GT10;
wire R18C34_GB70;
wire R1C47_X08;
wire R11C29_GBO0;
wire R28C31_SEL5;
wire R6C32_GB30;
wire R2C31_GBO1;
wire R28C28_N27;
wire R24C11_GBO1;
wire R5C33_GT00;
wire R10C25_E81;
wire R10C43_D2;
wire R28C7_E13;
wire R27C3_GB30;
wire R9C8_GB50;
wire R10C7_E27;
wire R25C39_GB50;
wire R5C39_GT00;
wire R17C37_GB20;
wire R28C19_E81;
wire R27C35_GB70;
wire R14C46_GB20;
wire R10C10_N80;
wire R10C40_E12;
wire R7C43_GT10;
wire R22C42_GB20;
wire R28C22_S23;
wire R10C26_C7;
wire R3C20_GB40;
wire R10C31_A4;
wire R10C10_LSR1;
wire R10C43_N23;
wire R10C43_B6;
wire R11C25_GT00;
wire R28C43_F2;
wire R10C29_UNK124;
wire R17C45_GT10;
wire R9C24_GB00;
wire R24C5_GB70;
wire R26C5_GB50;
wire R17C15_GB00;
wire R22C26_GB20;
wire R17C29_GB40;
wire R10C30_UNK126;
wire R4C20_GB00;
wire R4C8_GB50;
wire R10C43_C5;
wire R2C17_GB20;
wire R11C43_GBO1;
wire R21C43_GB60;
wire R10C16_D0;
wire R28C4_S82;
wire R6C14_GB10;
wire R28C25_F6;
wire R15C29_GB20;
wire R10C13_E27;
wire R8C44_GB00;
wire R4C11_GB50;
wire R17C22_GT00;
wire R26C15_GB70;
wire R10C19_SEL2;
wire R23C35_GB60;
wire R17C15_GT00;
wire R28C22_CE0;
wire R24C35_GB60;
wire R10C10_E27;
wire R8C27_GB10;
wire R13C2_GB10;
wire R17C38_GB10;
wire R12C43_GB20;
wire R10C40_W21;
wire R10C26_S24;
wire R10C27_X02;
wire R6C18_GB40;
wire R10C43_N25;
wire R5C32_GB00;
wire R23C18_GB40;
wire R24C4_GB00;
wire R10C34_W26;
wire R7C19_GB20;
wire R27C18_GB30;
wire R11C39_GBO1;
wire R23C33_GB60;
wire R20C5_GBO1;
wire R26C21_GB50;
wire R14C12_GB20;
wire R6C28_GB50;
wire R11C4_GT00;
wire R10C31_N20;
wire R21C32_GB70;
wire R28C31_D7;
wire R8C33_GB60;
wire R10C16_N10;
wire R12C22_GB50;
wire R27C39_GBO0;
wire R10C43_X02;
wire R29C28_C7;
wire R10C10_C0;
wire R21C28_GB00;
wire R4C32_GBO1;
wire R24C13_GB30;
wire R9C37_GB00;
wire R7C38_GB40;
wire R22C43_GB20;
wire R10C13_W82;
wire R12C7_GB70;
wire R10C34_A5;
wire R28C13_D1;
wire R10C31_Q6;
wire R28C28_S11;
wire R28C37_SEL3;
wire R10C22_W82;
wire R11C29_GB20;
wire R23C24_GT10;
wire R2C6_GT00;
wire R14C18_GB10;
wire R7C2_GB50;
wire R11C21_GT10;
wire R10C22_A3;
wire R9C23_GB40;
wire R8C24_GB60;
wire R6C27_GT10;
wire R1C47_N21;
wire R28C25_LSR2;
wire R10C34_F7;
wire R15C30_GB00;
wire R7C12_GB00;
wire R2C12_GT00;
wire R12C17_GT10;
wire R22C40_GBO0;
wire R28C10_SEL6;
wire R28C25_D1;
wire R28C28_F3;
wire R13C19_GB50;
wire R1C32_S81;
wire R10C26_N12;
wire R15C25_GBO0;
wire R1C47_SEL1;
wire R10C7_S26;
wire R28C4_X08;
wire R28C34_X06;
wire R10C16_S12;
wire R20C10_SPINE18;
wire R10C40_E82;
wire R4C29_GB40;
wire R14C40_GB00;
wire R28C40_F6;
wire R29C28_F1;
wire R25C37_GBO0;
wire R6C7_GT00;
wire R22C20_GB70;
wire R17C14_GBO0;
wire R1C28_W83;
wire R28C22_S24;
wire R6C39_GBO0;
wire R11C2_GB70;
wire R7C8_GBO0;
wire R20C18_GB50;
wire R10C25_N20;
wire R20C19_GB00;
wire R12C16_GT00;
wire R22C28_GB40;
wire R14C1_GT10;
wire R17C36_GBO0;
wire R10C31_S11;
wire R28C7_E82;
wire R8C10_GBO0;
wire R10C40_Q3;
wire R2C20_GBO1;
wire R22C45_GB10;
wire R17C38_GB30;
wire R1C47_S20;
wire R28C13_X03;
wire R18C13_GBO0;
wire R10C26_A5;
wire R26C16_GT10;
wire R5C8_GB70;
wire R17C29_GBO0;
wire R4C8_GB70;
wire R2C34_GBO1;
wire R24C23_GB10;
wire R10C27_W13;
wire R2C2_GT00;
wire R10C30_N12;
wire R13C20_GB70;
wire R28C22_F3;
wire R10C28_S20;
wire R28C34_A4;
wire R28C25_CE0;
wire R5C33_GB10;
wire R20C24_SPINE16;
wire R10C26_Q6;
wire R3C13_GB60;
wire R10C19_S21;
wire R10C19_E24;
wire R28C37_CLK2;
wire R24C33_GB20;
wire R24C29_GB30;
wire R27C37_GB10;
wire R21C18_GB50;
wire R7C37_GB50;
wire R14C11_GB60;
wire R13C18_GB50;
wire R2C1_SPINE11;
wire R22C36_GB30;
wire R3C30_GB30;
wire R3C11_GB10;
wire R15C38_GBO0;
wire R20C43_GB50;
wire R1C28_B7;
wire R10C13_B7;
wire R4C44_GBO0;
wire R10C19_E11;
wire R9C39_GBO1;
wire R24C3_GB60;
wire R1C1_N80;
wire R7C42_GT00;
wire R15C3_GB10;
wire R2C45_GT10;
wire R5C11_GB40;
wire R15C22_GBO1;
wire R14C11_GB50;
wire R3C29_GB60;
wire R13C31_GBO1;
wire R4C33_GBO1;
wire R10C13_D2;
wire R1C1_F3;
wire R10C16_W24;
wire R18C44_GB50;
wire R21C9_GT10;
wire R26C39_GBO0;
wire R28C22_S27;
wire R28C25_W12;
wire R28C40_D2;
wire R28C19_B7;
wire R20C22_GB30;
wire R28C7_LSR1;
wire R24C17_GB40;
wire R28C7_S22;
wire R28C28_D1;
wire R28C28_D6;
wire R26C35_GT10;
wire R18C14_GBO0;
wire R20C21_GBO0;
wire R26C6_GT10;
wire R18C21_GB50;
wire R1C1_W81;
wire R28C46_W80;
wire R1C32_S25;
wire R29C28_E80;
wire R10C19_N13;
wire R4C35_GT10;
wire R20C8_GB60;
wire R10C10_Q0;
wire R10C37_A2;
wire R24C23_GB50;
wire R28C46_E20;
wire R6C42_GB70;
wire R18C30_GB00;
wire R18C27_GB10;
wire R10C10_SN20;
wire R28C13_D5;
wire R13C34_GT10;
wire R24C28_GB30;
wire R22C4_GB30;
wire R16C22_GB40;
wire R21C45_GBO0;
wire R21C38_GB50;
wire R1C32_N11;
wire R4C7_GB20;
wire R20C30_SPINE26;
wire R10C16_EW10;
wire R10C29_D7;
wire R28C19_W27;
wire R28C40_S20;
wire R18C16_GB00;
wire R27C31_GBO1;
wire R6C22_GB20;
wire R14C38_GB20;
wire R24C40_GB50;
wire R10C40_Q6;
wire R16C11_GBO1;
wire R24C14_GT00;
wire R23C15_GB60;
wire R24C32_GB70;
wire R22C40_GB60;
wire R10C7_X07;
wire R2C17_GB50;
wire R20C13_GBO0;
wire R10C37_E21;
wire R20C32_SPINE28;
wire R10C40_N83;
wire R3C45_GBO0;
wire R1C28_F3;
wire R18C34_GB10;
wire R26C38_GB40;
wire R10C27_N25;
wire R20C2_GB40;
wire R23C30_GB70;
wire R28C31_A2;
wire R17C27_GB20;
wire R28C13_C7;
wire R27C13_GB50;
wire R17C23_GT00;
wire R9C39_GB50;
wire R20C13_GB60;
wire R5C3_GB60;
wire R15C29_GT10;
wire R11C7_GB60;
wire R18C8_GBO1;
wire R28C22_W21;
wire R28C43_C1;
wire R1C32_B2;
wire R7C35_GT00;
wire R20C20_GB70;
wire R28C43_EW10;
wire R28C28_S80;
wire R18C46_GB20;
wire R28C10_CLK0;
wire R15C30_GB10;
wire R21C9_GBO1;
wire R27C36_GBO1;
wire R17C22_GB40;
wire R20C22_GB50;
wire R18C9_GBO1;
wire R5C3_GT00;
wire R10C22_W13;
wire R25C14_GBO1;
wire R23C19_GB20;
wire R26C17_GB40;
wire R10C13_D6;
wire R6C36_GB10;
wire R17C26_GBO0;
wire R10C31_SEL3;
wire R14C34_GB50;
wire R26C5_GT00;
wire R11C44_GBO1;
wire R2C46_SPINE2;
wire R28C34_Q0;
wire R20C15_GB10;
wire R26C15_GBO0;
wire R9C5_GBO1;
wire R7C40_GB20;
wire R21C31_GB60;
wire R11C16_GBO1;
wire R6C17_GB40;
wire R10C37_Q5;
wire R25C13_GT10;
wire R6C8_GB70;
wire R25C9_GB10;
wire R3C15_GB40;
wire R10C27_C3;
wire R7C29_GB50;
wire R10C7_A4;
wire R18C34_GT10;
wire R10C30_W81;
wire R28C16_W12;
wire R28C31_CE0;
wire R16C5_GT00;
wire R20C13_GB40;
wire R17C41_GB10;
wire R28C19_X08;
wire R28C10_B6;
wire R5C25_GT00;
wire R25C6_GB00;
wire R26C7_GB10;
wire R2C20_GB10;
wire R27C43_GBO1;
wire R28C10_SEL1;
wire R17C19_GB20;
wire R23C9_GB20;
wire R3C26_GB60;
wire R8C42_GB00;
wire R15C20_GB40;
wire R10C37_B0;
wire R4C28_GB20;
wire R8C31_GB50;
wire R28C46_E82;
wire R7C45_GB70;
wire R27C39_GT10;
wire R21C22_GT10;
wire R14C33_GB00;
wire R1C32_W10;
wire R7C35_GB70;
wire R1C32_C0;
wire R6C12_GT10;
wire R21C25_GB10;
wire R12C42_GBO0;
wire R12C23_GB40;
wire R10C40_D4;
wire R26C32_GB70;
wire R20C44_GBO0;
wire R15C15_GT10;
wire R10C7_SEL3;
wire R2C14_GB60;
wire R22C5_GB20;
wire R20C26_GBO1;
wire R9C13_GB30;
wire R22C10_GBO0;
wire R26C40_GB70;
wire R8C26_GT00;
wire R9C5_GB20;
wire R6C32_GB40;
wire R20C8_SPINE16;
wire R13C27_GT00;
wire R2C45_GB10;
wire R20C32_GBO1;
wire R16C45_GB40;
wire R17C17_GT00;
wire R10C16_S27;
wire R23C5_GB50;
wire R3C43_GB10;
wire R20C35_GB20;
wire R21C45_GB10;
wire R26C9_GB50;
wire R5C37_GB00;
wire R10C13_E26;
wire R28C28_C7;
wire R21C4_GBO0;
wire R4C29_GB60;
wire R28C31_Q3;
wire R23C35_GB20;
wire R28C31_B6;
wire R28C4_SEL5;
wire R3C3_GB70;
wire R17C26_GB10;
wire R12C36_GB10;
wire R28C40_D4;
wire R1C47_EW20;
wire R20C12_GB60;
wire R7C21_GT10;
wire R22C23_GB50;
wire R3C20_GBO0;
wire R2C45_GBO0;
wire R22C7_GT10;
wire R27C40_GBO0;
wire R1C1_E81;
wire R23C16_GB00;
wire R10C30_C1;
wire R28C16_N82;
wire R2C27_GB70;
wire R25C2_GB20;
wire R23C45_GB30;
wire R2C11_GB40;
wire R23C27_GB60;
wire R13C24_GB30;
wire R17C11_GB00;
wire R24C40_GB20;
wire R10C7_Q5;
wire R21C1_GBO1;
wire R2C43_GB50;
wire R20C24_GT10;
wire R5C30_GB70;
wire R13C21_GB10;
wire R16C11_GB20;
wire R10C19_SN10;
wire R10C27_A1;
wire R6C25_GB20;
wire R26C46_GB00;
wire R10C34_C4;
wire R18C42_GB40;
wire R8C36_GBO1;
wire R10C30_CE1;
wire R28C25_CLK0;
wire R7C6_GB40;
wire R22C17_GB50;
wire R7C26_GB10;
wire R25C4_GBO0;
wire R16C21_GBO1;
wire R26C39_GB40;
wire R14C8_GB70;
wire R12C20_GBO0;
wire R21C42_GBO0;
wire R26C29_GB70;
wire R10C16_N23;
wire R3C45_GB10;
wire R9C26_GB70;
wire R8C11_GT10;
wire R7C12_GT00;
wire R28C31_D3;
wire R4C19_GB30;
wire R22C3_GT00;
wire R26C32_GT00;
wire R4C5_GB50;
wire R15C9_GB50;
wire R12C23_GB50;
wire R20C40_GB40;
wire R5C45_GB70;
wire R23C26_GB20;
wire R9C31_GT10;
wire R10C27_SN20;
wire R27C8_GBO0;
wire R1C28_S21;
wire R21C20_GB30;
wire R16C33_GB60;
wire R13C41_GB60;
wire R2C13_GT10;
wire R9C26_GB40;
wire R13C42_GB00;
wire R25C31_GBO1;
wire R24C30_GB50;
wire R21C37_GBO0;
wire R20C38_GBO1;
wire R10C31_CLK1;
wire R22C39_GB40;
wire R20C2_SPINE18;
wire R9C17_GT10;
wire R3C38_GBO1;
wire R17C46_GBO1;
wire R10C19_N24;
wire R18C11_GB60;
wire R4C20_GB70;
wire R18C34_GB30;
wire R6C39_GT10;
wire R1C1_W83;
wire R17C7_GT10;
wire R2C14_GBO0;
wire R10C22_W11;
wire R28C25_E81;
wire R16C40_GB50;
wire R14C2_GBO0;
wire R17C28_GB50;
wire R14C7_GB00;
wire R13C5_GB20;
wire R26C23_GB40;
wire R15C29_GB50;
wire R28C43_Q6;
wire R24C4_GB60;
wire R10C43_X07;
wire R28C16_S81;
wire R16C41_GBO1;
wire R28C43_D1;
wire R22C32_GB00;
wire R4C7_GB50;
wire R11C45_GB40;
wire R26C45_GB20;
wire R28C34_B7;
wire R3C21_GB30;
wire R16C3_GB50;
wire R6C33_GT00;
wire R12C45_GT10;
wire R27C45_GT00;
wire R11C46_GBO1;
wire R28C7_B4;
wire R1C47_A7;
wire R16C30_GB20;
wire R8C30_GBO1;
wire R14C9_GB70;
wire R13C16_GT10;
wire R21C12_GB20;
wire R13C33_GB00;
wire R28C43_F7;
wire R11C44_GB30;
wire R14C37_GB00;
wire R28C31_N13;
wire R14C26_GB30;
wire R16C12_GB70;
wire R20C26_GB30;
wire R21C13_GBO1;
wire R2C8_GBO0;
wire R10C7_B5;
wire R6C11_GB10;
wire R11C34_GB60;
wire R10C30_F3;
wire R10C26_A3;
wire R21C5_GB50;
wire R9C20_GBO0;
wire R25C41_GBO1;
wire R28C37_E20;
wire R26C30_GT10;
wire R10C22_N12;
wire R10C13_W21;
wire R12C21_GB00;
wire R25C41_GB10;
wire R24C19_GB40;
wire R12C33_GB20;
wire R8C7_GT00;
wire R8C30_GB70;
wire R2C40_GB70;
wire R10C22_N13;
wire R7C45_GBO0;
wire R16C42_GB00;
wire R10C30_C7;
wire R23C14_GB30;
wire R18C9_GB60;
wire R18C31_GBO0;
wire R7C38_GB50;
wire R13C38_GB60;
wire R28C25_E26;
wire R28C22_S82;
wire R18C38_GB50;
wire R20C45_GB60;
wire R9C21_GB00;
wire R28C31_SN20;
wire R2C7_GB60;
wire R28C46_EW10;
wire R7C5_GB20;
wire R10C28_E21;
wire R6C4_GB10;
wire R5C13_GT00;
wire R12C22_GT10;
wire R2C1_GBO1;
wire R11C34_GB70;
wire R1C32_W22;
wire R3C34_GB50;
wire R5C41_GB00;
wire R10C43_CE2;
wire R5C41_GB70;
wire R18C46_GT00;
wire R9C9_GT10;
wire R20C32_GT00;
wire R23C18_GB00;
wire R18C31_GB50;
wire R5C25_GB60;
wire R8C45_GB60;
wire R13C3_GB30;
wire R6C5_GT00;
wire R21C22_GB50;
wire R5C10_GB10;
wire R21C42_GT10;
wire R20C36_GB30;
wire R18C10_GT00;
wire R10C19_C0;
wire R10C40_W23;
wire R10C29_SEL4;
wire R21C32_GBO1;
wire R17C35_GBO1;
wire R10C29_B6;
wire R28C43_W82;
wire R28C28_W12;
wire R4C18_GB00;
wire R23C10_GBO1;
wire R16C18_GB00;
wire R10C34_E21;
wire R28C13_N11;
wire R5C6_GBO0;
wire R28C37_SN10;
wire R4C23_GB40;
wire R21C16_GT00;
wire R16C46_GBO1;
wire R8C22_GB30;
wire R12C44_GBO1;
wire R2C16_GB60;
wire R4C15_GT10;
wire R8C16_GB00;
wire R4C16_GT00;
wire R4C22_GBO0;
wire R6C12_GB30;
wire R11C4_GB00;
wire R4C34_GB30;
wire R6C31_GT10;
wire R25C23_GB50;
wire R12C36_GBO1;
wire R27C30_GBO0;
wire R1C28_LSR0;
wire R28C40_N82;
wire R10C27_D7;
wire R16C2_GB70;
wire R24C14_GB50;
wire R2C39_GB50;
wire R9C15_GBO1;
wire R28C16_LSR0;
wire R10C31_N11;
wire R5C27_GB10;
wire R27C32_GBO1;
wire R25C35_GB30;
wire R12C44_GT10;
wire R28C34_D2;
wire R22C6_GB30;
wire R3C43_GB30;
wire R27C24_GB30;
wire R3C45_GT00;
wire R20C31_SPINE25;
wire R9C16_GT10;
wire R5C20_GBO0;
wire R21C33_GT00;
wire R3C2_GB70;
wire R8C32_GB40;
wire R13C45_GB00;
wire R26C36_GB20;
wire R11C18_GB20;
wire R24C44_GB20;
wire R4C20_GBO0;
wire R18C9_GT10;
wire R4C33_GB30;
wire R12C31_GB20;
wire R25C37_GT00;
wire R16C42_GB20;
wire R2C4_GB20;
wire R10C19_B0;
wire R2C23_GB00;
wire R21C41_GB70;
wire R22C24_GT10;
wire R2C2_GB50;
wire R22C31_GB70;
wire R10C22_N21;
wire R3C22_GB60;
wire R5C3_GB50;
wire R28C16_B4;
wire R2C42_SPINE2;
wire R26C22_GB10;
wire R14C25_GB40;
wire R27C39_GB10;
wire R3C46_GBO1;
wire R7C30_GT10;
wire R21C2_GB40;
wire R3C44_GB60;
wire R28C16_E80;
wire R7C23_GBO0;
wire R15C18_GBO0;
wire R16C33_GB20;
wire R20C36_GB70;
wire R28C43_S22;
wire R23C41_GB60;
wire R3C9_GB40;
wire R1C1_S10;
wire R28C16_A3;
wire R28C43_F4;
wire R2C8_GB50;
wire R9C29_GT00;
wire R11C8_GT10;
wire R12C17_GBO0;
wire R12C12_GB30;
wire R8C29_GB50;
wire R7C19_GB30;
wire R14C3_GT00;
wire R5C29_GBO0;
wire R17C19_GB60;
wire R8C42_GB30;
wire R18C19_GB50;
wire R1C28_A5;
wire R28C40_C4;
wire R28C31_LSR0;
wire R1C1_N21;
wire R2C13_GT00;
wire R6C39_GB10;
wire R11C25_GB70;
wire R10C34_E12;
wire R8C5_GB30;
wire R1C1_X04;
wire R3C22_GB20;
wire R10C16_E20;
wire R14C20_GB30;
wire R26C7_GB40;
wire R21C21_GB10;
wire R7C41_GBO1;
wire R18C43_GB20;
wire R20C2_GBO1;
wire R2C28_GB00;
wire R16C13_GB40;
wire R28C43_E81;
wire R8C37_GBO1;
wire R28C43_Q4;
wire R6C8_GB50;
wire R2C25_GT10;
wire R11C31_GBO1;
wire R20C46_GB00;
wire R21C37_GB50;
wire R6C27_GB70;
wire R15C10_GT00;
wire R24C39_GB70;
wire R28C7_D5;
wire R9C26_GT00;
wire R2C27_GBO1;
wire R10C13_A2;
wire R9C22_GBO1;
wire R10C29_SEL7;
wire R24C25_GB10;
wire R12C30_GB20;
wire R10C31_EW20;
wire R11C29_GB60;
wire R2C26_GB10;
wire R13C7_GB00;
wire R21C32_GB50;
wire R11C17_GB70;
wire R15C40_GB70;
wire R9C34_GT10;
wire R13C11_GT10;
wire R21C29_GT00;
wire R3C37_GBO1;
wire R7C22_GB10;
wire R10C28_CE0;
wire R15C16_GB40;
wire R1C47_F3;
wire R7C46_GB50;
wire R10C10_N81;
wire R6C29_GT00;
wire R10C22_E13;
wire R3C29_GB30;
wire R13C40_GBO0;
wire R20C42_SPINE26;
wire R28C28_B4;
wire R20C18_GBO1;
wire R17C10_GB20;
wire R16C38_GB30;
wire R2C25_GBO0;
wire R15C18_GB60;
wire R25C36_GBO0;
wire R27C2_GB30;
wire R10C16_Q2;
wire R13C5_GB50;
wire R22C44_GBO0;
wire R7C22_GB50;
wire R29C28_C0;
wire R23C19_GT10;
wire R15C7_GT00;
wire R20C31_GB20;
wire R11C41_GB20;
wire R10C43_SEL7;
wire R10C29_E80;
wire R7C3_GB60;
wire R27C9_GB20;
wire R16C18_GB70;
wire R17C19_GB40;
wire R10C27_W81;
wire R4C37_GB40;
wire R28C7_B6;
wire R14C45_GB10;
wire R10C43_E27;
wire R4C25_GBO1;
wire R7C15_GB30;
wire R7C45_GBO1;
wire R20C6_GT00;
wire R24C29_GB70;
wire R13C46_GB70;
wire R28C46_SEL5;
wire R1C47_E21;
wire R13C21_GB50;
wire R20C18_GB30;
wire R7C43_GB00;
wire R18C36_GB10;
wire R1C32_CLK2;
wire R10C29_F6;
wire R25C11_GBO0;
wire R16C5_GB70;
wire R28C19_Q3;
wire R28C10_Q7;
wire R12C38_GB30;
wire R14C42_GB10;
wire R26C6_GBO0;
wire R28C16_N25;
wire R1C47_S23;
wire R28C31_N12;
wire R24C5_GB60;
wire R7C23_GB10;
wire R20C26_GB00;
wire R22C41_GB30;
wire R17C32_GB40;
wire R1C47_SEL4;
wire R10C7_A6;
wire R15C16_GBO0;
wire R28C10_D5;
wire R21C4_GB60;
wire R5C6_GB10;
wire R4C41_GB20;
wire R22C9_GT10;
wire R10C31_E80;
wire R10C10_N83;
wire R10C25_W24;
wire R28C40_EW20;
wire R21C34_GT00;
wire R28C16_S12;
wire R5C15_GB20;
wire R8C29_GBO0;
wire R17C17_GT10;
wire R24C3_GB40;
wire R26C2_GB70;
wire R3C35_GB70;
wire R22C43_GB70;
wire R24C6_GB50;
wire R28C16_Q6;
wire R1C32_W21;
wire R4C42_GB50;
wire R28C34_D1;
wire R16C23_GB20;
wire R28C37_E80;
wire R14C45_GB70;
wire R11C5_GBO0;
wire R21C43_GT10;
wire R8C13_GB00;
wire R18C35_GBO0;
wire R16C9_GB40;
wire R1C32_N21;
wire R26C26_GBO1;
wire R8C9_GT10;
wire R28C43_C0;
wire R8C46_GB30;
wire R9C3_GB60;
wire R28C28_C6;
wire R14C32_GB70;
wire R23C11_GB50;
wire R26C14_GB50;
wire R27C21_GB70;
wire R27C4_GB60;
wire R22C41_GB00;
wire R28C34_E23;
wire R28C19_W82;
wire R7C5_GT10;
wire R28C10_S83;
wire R28C31_C1;
wire R5C10_GB40;
wire R12C3_GB20;
wire R10C19_E13;
wire R10C34_W82;
wire R14C30_GB60;
wire R12C31_GB10;
wire R10C10_S27;
wire R5C5_GB70;
wire R10C34_C7;
wire R22C35_GT00;
wire R10C28_LSR0;
wire R28C40_N10;
wire R11C35_GBO1;
wire R5C28_GB00;
wire R18C25_GB30;
wire R27C46_GB50;
wire R10C27_CE2;
wire R10C34_Q0;
wire R8C7_GB10;
wire R28C46_E80;
wire R21C34_GB60;
wire R8C14_GB10;
wire R28C25_X08;
wire R24C11_GB70;
wire R13C5_GB30;
wire R13C16_GB20;
wire R9C33_GB40;
wire R29C28_A1;
wire R14C26_GB40;
wire R10C16_C3;
wire R9C39_GB40;
wire R4C5_GB40;
wire R2C29_GB30;
wire R28C37_CE1;
wire R8C15_GT00;
wire R8C38_GT00;
wire R17C39_GB30;
wire R6C3_GB70;
wire R3C44_GB00;
wire R1C28_X01;
wire R28C43_X05;
wire R24C20_GB70;
wire R5C41_GB30;
wire R2C44_GB40;
wire R4C15_GT00;
wire R8C16_GB60;
wire R10C16_C0;
wire R3C7_GBO1;
wire R21C5_GB30;
wire R5C31_GB00;
wire R27C43_GB20;
wire R10C37_N22;
wire R7C31_GB30;
wire R23C33_GB20;
wire R24C8_GB40;
wire R15C45_GT00;
wire R10C28_Q5;
wire R24C26_GB70;
wire R14C5_GBO0;
wire R12C29_GB20;
wire R26C21_GB20;
wire R20C28_GB70;
wire R6C26_GB30;
wire R18C26_GT00;
wire R10C7_C0;
wire R2C5_GBO1;
wire R27C2_GBO1;
wire R14C34_GB40;
wire R26C43_GB70;
wire R10C10_SEL7;
wire R17C31_GB70;
wire R12C12_GT00;
wire R10C40_E21;
wire R1C32_B1;
wire R22C34_GB00;
wire R28C40_W11;
wire R23C39_GB40;
wire R13C9_GB30;
wire R16C10_GB40;
wire R24C26_GB50;
wire R6C27_GB60;
wire R17C38_GBO1;
wire R28C43_N10;
wire R10C10_CE2;
wire R20C24_GB70;
wire R9C30_GBO1;
wire R16C39_GT10;
wire R10C22_S21;
wire R24C41_GB10;
wire R8C2_GB60;
wire R11C10_GBO1;
wire R10C26_S82;
wire R24C15_GB30;
wire R13C23_GT00;
wire R17C4_GB60;
wire R26C5_GBO1;
wire R27C37_GB30;
wire R1C1_E26;
wire R23C14_GBO0;
wire R10C10_A0;
wire R28C28_N22;
wire R28C10_B7;
wire R28C7_X03;
wire R9C46_GB20;
wire R24C41_GB00;
wire R10C43_SEL4;
wire R28C16_SEL6;
wire R4C16_GBO0;
wire R9C19_GB70;
wire R7C36_GB30;
wire R15C7_GT10;
wire R4C36_GB60;
wire R28C7_W24;
wire R6C39_GB70;
wire R3C34_GBO1;
wire R7C43_GB40;
wire R8C18_GB60;
wire R7C41_GBO0;
wire R25C41_GB30;
wire R26C34_GBO1;
wire R22C11_GB70;
wire R3C35_GB00;
wire R15C33_GB70;
wire R28C28_EW20;
wire R10C25_W80;
wire R2C3_GT10;
wire R21C25_GB70;
wire R4C38_GB10;
wire R2C36_GB20;
wire R14C40_GB70;
wire R10C26_W27;
wire R13C29_GB30;
wire R10C10_W24;
wire R10C31_S20;
wire R18C35_GT10;
wire R20C1_GT00;
wire R14C22_GBO1;
wire R21C31_GB50;
wire R2C19_GB40;
wire R10C13_N81;
wire R8C37_GB40;
wire R28C16_EW10;
wire R15C3_GB40;
wire R15C31_GB40;
wire R25C24_GBO0;
wire R5C34_GB20;
wire R20C5_GB00;
wire R10C7_W80;
wire R13C36_GT00;
wire R11C7_GB50;
wire R17C30_GB20;
wire R9C8_GB40;
wire R29C29_F6;
wire R25C15_GB70;
wire R5C7_GB40;
wire R20C35_GBO1;
wire R1C47_N80;
wire R3C8_GB00;
wire R24C10_GB60;
wire R6C28_GB10;
wire R13C32_GB40;
wire R25C19_GT00;
wire R25C34_GB50;
wire R10C30_B3;
wire R5C11_GB20;
wire R11C29_GT00;
wire R23C12_GB30;
wire R16C38_GB20;
wire R1C28_B3;
wire R28C25_X01;
wire R15C28_GB50;
wire R4C8_GB40;
wire R28C25_B4;
wire R14C3_GBO1;
wire R10C7_X08;
wire R24C36_GB30;
wire R20C36_GBO1;
wire R10C37_E27;
wire R3C1_GBO0;
wire R17C44_GT10;
wire R21C27_GB00;
wire R5C44_GB40;
wire R10C40_S25;
wire R27C35_GB40;
wire R23C35_GBO1;
wire R22C36_GT10;
wire R24C6_GB70;
wire R27C43_GB60;
wire R14C37_GB70;
wire R18C14_GB50;
wire R15C37_GB60;
wire R28C16_LSR1;
wire R8C5_GB10;
wire R16C13_GB30;
wire R26C25_GB50;
wire R8C42_GB40;
wire R10C16_X03;
wire R16C22_GBO1;
wire R10C29_SEL5;
wire R27C5_GB00;
wire R10C27_UNK121;
wire R28C31_CE2;
wire R15C12_GB30;
wire R11C41_GBO1;
wire R12C41_GB10;
wire R11C4_GB10;
wire R12C16_GB20;
wire R9C10_GB20;
wire R7C4_GB60;
wire R26C18_GBO1;
wire R16C31_GBO1;
wire R28C40_X07;
wire R2C18_GB50;
wire R7C14_GB30;
wire R22C23_GB40;
wire R28C34_W83;
wire R22C1_GT10;
wire R28C22_CE2;
wire R4C26_GB60;
wire R22C19_GB20;
wire R12C10_GB70;
wire R13C15_GB30;
wire R6C29_GB60;
wire R4C36_GB70;
wire R5C11_GB00;
wire R22C34_GB20;
wire R12C39_GB30;
wire R3C27_GT00;
wire R2C33_GB30;
wire R20C38_GB40;
wire R15C8_GT00;
wire R11C35_GT10;
wire R11C15_GB10;
wire R5C3_GB20;
wire R27C24_GB00;
wire R27C3_GBO0;
wire R11C24_GB50;
wire R14C41_GB70;
wire R8C40_GB00;
wire R1C1_E25;
wire R28C16_S23;
wire R22C15_GB70;
wire R27C1_GBO0;
wire R10C13_SEL6;
wire R13C41_GT10;
wire R28C4_W12;
wire R3C37_GT10;
wire R13C13_GB20;
wire R20C12_GBO1;
wire R26C2_GT00;
wire R14C14_GB70;
wire R4C35_GB20;
wire R10C29_CLK2;
wire R9C8_GBO0;
wire R28C34_X07;
wire R8C2_GT10;
wire R17C28_GB40;
wire R29C28_SEL1;
wire R26C3_GB20;
wire R11C21_GB20;
wire R3C38_GB50;
wire R26C44_GBO0;
wire R17C5_GB40;
wire R26C37_GB70;
wire R15C9_GT00;
wire R28C40_N24;
wire R26C28_GB20;
wire R15C46_GB30;
wire R29C28_N11;
wire R5C35_GB70;
wire R28C37_E21;
wire R17C33_GB20;
wire R9C18_GT10;
wire R2C30_GB30;
wire R17C31_GT10;
wire R24C1_GT10;
wire R29C28_Q2;
wire R3C2_GB30;
wire R10C28_CE2;
wire R25C11_GB50;
wire R15C20_GT00;
wire R4C38_GT10;
wire R10C7_W25;
wire R8C28_GB50;
wire R7C31_GT00;
wire R6C43_GB40;
wire R10C31_B2;
wire R10C19_S11;
wire R26C15_GBO1;
wire R8C14_GB70;
wire R27C5_GB20;
wire R13C44_GB20;
wire R15C45_GBO0;
wire R10C28_F2;
wire R15C5_GBO0;
wire R26C23_GB60;
wire R12C26_GB60;
wire R23C30_GB20;
wire R1C32_W12;
wire R10C43_D4;
wire R28C40_N25;
wire R4C43_GT00;
wire R17C7_GB20;
wire R12C20_GB30;
wire R11C15_GB50;
wire R4C2_GB30;
wire R7C11_GB30;
wire R26C4_GB60;
wire R1C47_D4;
wire R14C23_GB10;
wire R28C43_F1;
wire R26C23_GB20;
wire R16C6_GB30;
wire R26C46_GB10;
wire R10C13_E20;
wire R28C40_A2;
wire R14C26_GT00;
wire R4C33_GT10;
wire R16C26_GB70;
wire R10C31_F3;
wire R22C25_GBO1;
wire R13C17_GB20;
wire R21C19_GB70;
wire R13C38_GB00;
wire R14C46_GB10;
wire R25C36_GT10;
wire R22C39_GBO1;
wire R10C22_EW10;
wire R21C45_GB50;
wire R28C31_A3;
wire R18C28_GB70;
wire R6C45_GB40;
wire R25C25_GB20;
wire R6C32_GBO0;
wire R17C45_GB60;
wire R15C27_GB60;
wire R27C27_GB10;
wire R8C12_GB60;
wire R7C9_GB30;
wire R3C10_GB40;
wire R5C26_GB70;
wire R10C7_S20;
wire R4C45_GT10;
wire R28C7_CLK1;
wire R17C29_GB60;
wire R8C17_GBO0;
wire R28C40_W83;
wire R10C29_X01;
wire R16C32_GB00;
wire R21C24_GB40;
wire R28C10_C3;
wire R8C2_GT00;
wire R15C44_GB00;
wire R3C30_GT00;
wire R7C37_GBO0;
wire R10C26_E81;
wire R10C43_E10;
wire R5C27_GT00;
wire R28C7_B1;
wire R3C5_GB20;
wire R24C12_GB00;
wire R23C32_GB00;
wire R2C7_GB00;
wire R18C45_GT00;
wire R12C16_GB40;
wire R5C17_GB50;
wire R3C38_GT00;
wire R26C14_GB30;
wire R17C43_GB40;
wire R28C40_X02;
wire R18C21_GT10;
wire R9C36_GT00;
wire R4C14_GBO1;
wire R1C47_E82;
wire R10C22_C4;
wire R2C10_GB60;
wire R18C33_GB50;
wire R12C42_GB00;
wire R10C19_B6;
wire R13C28_GB30;
wire R17C46_GT00;
wire R25C9_GBO1;
wire R11C24_GT10;
wire R17C23_GBO1;
wire R23C34_GBO0;
wire R16C44_GBO0;
wire R10C13_A6;
wire R13C18_GB60;
wire R14C26_GB60;
wire R5C41_GB60;
wire R10C16_N22;
wire R11C12_GB20;
wire R11C5_GB50;
wire R10C43_N80;
wire R6C15_GB00;
wire R23C17_GB40;
wire R7C12_GB10;
wire R5C27_GB00;
wire R6C41_GB60;
wire R24C18_GB50;
wire R9C2_GBO1;
wire R1C47_S24;
wire R28C10_E22;
wire R2C46_GB70;
wire R26C43_GB40;
wire R10C16_D7;
wire R2C17_GB30;
wire R24C18_GT10;
wire R8C5_GB40;
wire R8C6_GT00;
wire R14C4_GB50;
wire R8C26_GB50;
wire R27C17_GBO0;
wire R14C24_GT10;
wire R24C18_GB30;
wire R23C42_GT00;
wire R7C15_GBO0;
wire R5C17_GB40;
wire R27C39_GB30;
wire R16C26_GBO1;
wire R12C24_GT10;
wire R11C8_GB40;
wire R6C40_GB40;
wire R28C4_B7;
wire R22C10_GB70;
wire R28C37_W13;
wire R1C32_SEL5;
wire R15C34_GB00;
wire R20C19_GBO1;
wire R25C35_GBO0;
wire R10C26_Q0;
wire R14C31_GB20;
wire R12C25_GB40;
wire R7C5_GBO0;
wire R25C42_GB40;
wire R7C45_GT00;
wire R6C43_GB00;
wire R1C28_Q6;
wire R4C10_GB00;
wire R24C30_GB00;
wire R6C3_GB50;
wire R23C30_GB60;
wire R5C28_GB70;
wire R26C15_GB30;
wire R13C28_GB70;
wire R25C28_GT00;
wire R26C42_GT00;
wire R28C37_E11;
wire R27C3_GB20;
wire R20C33_GB20;
wire R23C3_GB60;
wire R9C43_GT10;
wire R13C25_GB10;
wire R9C25_GB70;
wire R10C13_C4;
wire R28C7_EW10;
wire R28C22_S26;
wire R22C20_GB10;
wire R5C21_GB00;
wire R21C8_GB30;
wire R23C10_GB20;
wire R10C31_N22;
wire R13C24_GBO0;
wire R16C27_GBO1;
wire R10C31_E10;
wire R23C43_GB30;
wire R28C4_S10;
wire R18C3_GB10;
wire R25C34_GB10;
wire R28C31_W21;
wire R20C43_GBO0;
wire R9C28_GT10;
wire R13C2_GB70;
wire R1C28_N22;
wire R10C22_W23;
wire R10C31_SEL4;
wire R17C5_GB70;
wire R13C46_GB60;
wire R8C8_GT00;
wire R12C4_GT10;
wire R4C24_GB20;
wire R7C27_GB20;
wire R3C16_GB20;
wire R4C18_GBO0;
wire R8C23_GT00;
wire R22C1_GBO0;
wire R25C6_GB20;
wire R10C19_E22;
wire R10C19_W21;
wire R1C1_N81;
wire R28C34_A6;
wire R21C8_GB00;
wire R15C2_GT00;
wire R16C10_GB20;
wire R1C32_X04;
wire R28C37_C6;
wire R28C13_N83;
wire R20C22_SPINE18;
wire R5C14_GBO0;
wire R10C13_A4;
wire R10C43_S10;
wire R25C38_GBO1;
wire R20C41_GT10;
wire R7C29_GB60;
wire R1C47_E24;
wire R5C23_GB30;
wire R22C14_GB10;
wire R3C3_GBO0;
wire R10C26_W80;
wire R10C34_C3;
wire R14C30_GB50;
wire R11C38_GB60;
wire R25C21_GB10;
wire R4C16_GB50;
wire R10C29_Q7;
wire R7C31_GB60;
wire R25C39_GB70;
wire R2C44_GB10;
wire R17C39_GBO0;
wire R17C23_GB20;
wire R15C37_GT10;
wire R7C13_GB60;
wire R10C28_N11;
wire R10C37_S26;
wire R3C32_GT10;
wire R16C15_GB40;
wire R28C37_SEL6;
wire R8C38_GB60;
wire R13C11_GBO1;
wire R24C21_GB20;
wire R8C6_GB20;
wire R3C39_GB00;
wire R28C19_A4;
wire R17C5_GT00;
wire R21C41_GB30;
wire R21C20_GB40;
wire R21C45_GBO1;
wire R23C22_GB00;
wire R5C28_GB20;
wire R24C26_GB40;
wire R1C32_W82;
wire R27C2_GB10;
wire R28C16_SEL2;
wire R28C19_S23;
wire R28C40_X04;
wire R10C40_N13;
wire R7C13_GB20;
wire R18C8_GB60;
wire R4C19_GBO1;
wire R2C44_GB50;
wire R10C40_SEL6;
wire R10C29_W27;
wire R23C14_GT00;
wire R10C25_SEL6;
wire R18C4_GB50;
wire R17C19_GB50;
wire R16C22_GT10;
wire R6C4_GBO0;
wire R28C22_A3;
wire R6C16_GB10;
wire R14C14_GBO1;
wire R26C5_GT10;
wire R16C34_GB10;
wire R8C11_GB60;
wire R21C46_GB30;
wire R28C34_EW20;
wire R18C8_GT10;
wire R6C41_GBO1;
wire R20C43_SPINE29;
wire R26C26_GBO0;
wire R16C16_GB50;
wire R1C1_E83;
wire R1C28_SEL5;
wire R10C19_S24;
wire R22C39_GB50;
wire R28C19_S83;
wire R10C16_W27;
wire R28C7_C0;
wire R16C44_GBO1;
wire R28C34_SEL7;
wire R5C24_GB30;
wire R28C4_W23;
wire R11C17_GB00;
wire R1C47_Q7;
wire R10C28_D0;
wire R8C46_GBO1;
wire R2C13_GB60;
wire R26C33_GT10;
wire R3C14_GB00;
wire R4C12_GB00;
wire R9C20_GT10;
wire R5C15_GB40;
wire R10C26_N13;
wire R12C43_GB40;
wire R16C25_GB20;
wire R10C13_N13;
wire R10C26_CE1;
wire R28C16_A1;
wire R2C28_GT10;
wire R6C15_GB50;
wire R12C28_GT10;
wire R10C16_E23;
wire R11C5_GB20;
wire R16C28_GB60;
wire R3C33_GB30;
wire R23C13_GB70;
wire R8C10_GT10;
wire R23C10_GB00;
wire R11C41_GB10;
wire R13C21_GT00;
wire R10C43_F5;
wire R15C27_GBO1;
wire R11C27_GB30;
wire R28C31_X01;
wire R7C39_GBO1;
wire R1C32_W80;
wire R8C40_GB20;
wire R17C6_GB60;
wire R28C25_S27;
wire R6C40_GT00;
wire R13C41_GBO0;
wire R28C13_X04;
wire R24C11_GB50;
wire R26C38_GB10;
wire R28C4_C3;
wire R10C43_SN20;
wire R28C43_SEL5;
wire R10C10_N21;
wire R3C14_GB30;
wire R11C41_GB00;
wire R9C42_GT00;
wire R22C4_GB00;
wire R28C43_F6;
wire R22C20_GB60;
wire R14C24_GBO1;
wire R7C39_GT10;
wire R26C43_GBO0;
wire R10C34_E10;
wire R21C14_GB00;
wire R3C36_GB40;
wire R29C28_S24;
wire R28C43_B3;
wire R14C21_GB00;
wire R8C26_GB70;
wire R28C7_S26;
wire R2C7_GB70;
wire R9C37_GBO0;
wire R13C34_GB70;
wire R10C22_SEL7;
wire R10C29_F1;
wire R21C41_GT00;
wire R20C27_GB10;
wire R20C25_GB10;
wire R10C19_X03;
wire R21C9_GB30;
wire R15C20_GB20;
wire R10C34_A0;
wire R20C16_GBO0;
wire R7C8_GB30;
wire R6C23_GT10;
wire R25C26_GBO1;
wire R20C19_GBO0;
wire R11C33_GB00;
wire R23C46_GB50;
wire R28C31_E21;
wire R5C35_GBO0;
wire R28C19_A2;
wire R28C16_W27;
wire R17C12_GBO0;
wire R17C43_GB20;
wire R15C43_GB40;
wire R16C34_GT10;
wire R8C9_GB00;
wire R22C22_GB10;
wire R12C15_GB60;
wire R9C45_GB30;
wire R10C43_N22;
wire R26C31_GB00;
wire R1C28_S27;
wire R23C3_GB10;
wire R5C33_GB50;
wire R28C19_C1;
wire R11C20_GB70;
wire R10C43_SEL6;
wire R3C39_GB60;
wire R18C32_GB50;
wire R1C1_N10;
wire R13C43_GB10;
wire R12C23_GB70;
wire R10C19_Q4;
wire R10C31_SEL7;
wire R28C34_Q5;
wire R4C39_GB50;
wire R27C2_GT00;
wire R22C12_GB30;
wire R28C34_E81;
wire R10C37_N12;
wire R28C4_S83;
wire R11C33_GT10;
wire R10C13_N12;
wire R10C19_A6;
wire R3C2_GBO0;
wire R28C28_C2;
wire R18C3_GB20;
wire R3C35_GB40;
wire R28C40_W22;
wire R7C33_GT10;
wire R20C21_GB30;
wire R17C3_GB40;
wire R26C8_GB60;
wire R21C4_GB50;
wire R16C6_GB70;
wire R25C15_GB50;
wire R25C32_GBO1;
wire R28C4_W27;
wire R26C24_GB40;
wire R14C33_GBO0;
wire R14C27_GB50;
wire R28C31_S23;
wire R14C11_GBO1;
wire R9C32_GB40;
wire R2C28_GB10;
wire R7C3_GB30;
wire R5C10_GB50;
wire R26C17_GB60;
wire R24C6_GB40;
wire R23C36_GB20;
wire R10C16_CE1;
wire R1C32_A3;
wire R23C22_GB60;
wire R20C3_GB70;
wire R11C19_GB40;
wire R21C22_GT00;
wire R2C39_GB00;
wire R17C40_GT10;
wire R10C16_S83;
wire R10C26_C3;
wire R6C30_GBO1;
wire R6C46_GB70;
wire R14C4_GB40;
wire R10C16_F0;
wire R28C37_X01;
wire R11C30_GB70;
wire R21C6_GB20;
wire R10C27_E26;
wire R26C1_GT00;
wire R13C26_GB00;
wire R6C23_GB50;
wire R13C24_GB00;
wire R3C23_GB10;
wire R12C17_GB60;
wire R27C35_GBO0;
wire R1C28_W27;
wire R28C43_W13;
wire R26C6_GB60;
wire R21C32_GT10;
wire R8C39_GB60;
wire R24C22_GB30;
wire R23C44_GB30;
wire R28C10_Q3;
wire R22C39_GB10;
wire R9C21_GB20;
wire R2C6_GB30;
wire R17C46_GB00;
wire R10C25_F3;
wire R28C43_CLK0;
wire R28C34_B4;
wire R7C13_GB30;
wire R28C19_N82;
wire R13C32_GBO1;
wire R8C40_GBO1;
wire R2C27_GB40;
wire R12C38_GBO0;
wire R10C43_C7;
wire R10C19_N81;
wire R25C14_GB70;
wire R28C16_S83;
wire R14C20_GBO1;
wire R10C25_E83;
wire R20C40_GB00;
wire R13C31_GT10;
wire R25C14_GB10;
wire R13C14_GB30;
wire R5C16_GB00;
wire R7C24_GB10;
wire R10C16_N27;
wire R26C22_GT10;
wire R28C40_X03;
wire R23C14_GT10;
wire R26C19_GB50;
wire R4C18_GT10;
wire R10C37_A7;
wire R6C11_GB00;
wire R7C42_GB30;
wire R14C15_GT00;
wire R9C40_GB50;
wire R17C4_GB00;
wire R24C34_GT10;
wire R1C28_LSR2;
wire R5C14_GT00;
wire R5C26_GT10;
wire R26C27_GB60;
wire R20C39_GB10;
wire R25C11_GB40;
wire R6C14_GB40;
wire R8C8_GB50;
wire R26C18_GB20;
wire R15C38_GB10;
wire R7C38_GT10;
wire R22C5_GBO1;
wire R5C38_GBO0;
wire R5C3_GB30;
wire R7C36_GB10;
wire R18C4_GB10;
wire R6C46_GT10;
wire R25C45_GB50;
wire R10C40_N10;
wire R24C1_GT00;
wire R3C42_GB20;
wire R2C27_SPINE13;
wire R2C10_GB40;
wire R6C4_GB60;
wire R23C37_GB30;
wire R8C41_GT10;
wire R28C7_CE1;
wire R5C44_GT00;
wire R2C21_GB30;
wire R8C40_GB60;
wire R8C4_GB60;
wire R8C44_GB20;
wire R1C32_C3;
wire R3C5_GBO1;
wire R9C15_GB60;
wire R15C14_GB10;
wire R10C28_W27;
wire R10C26_X04;
wire R10C27_UNK124;
wire R27C38_GB60;
wire R28C34_F3;
wire R28C4_E21;
wire R6C34_GBO1;
wire R10C37_N26;
wire R10C27_SPINE12;
wire R28C25_N13;
wire R4C20_GB10;
wire R3C23_GBO0;
wire R16C24_GT00;
wire R9C2_GB30;
wire R1C1_CLK2;
wire R7C23_GB50;
wire R9C43_GB10;
wire R7C25_GB10;
wire R12C11_GBO0;
wire R25C11_GB20;
wire R26C4_GB00;
wire R7C22_GB30;
wire R23C28_GB10;
wire R27C11_GB30;
wire R28C31_N81;
wire R27C25_GB00;
wire R28C40_SEL3;
wire R29C28_E21;
wire R10C10_CLK2;
wire R28C34_W20;
wire R24C46_GBO0;
wire R22C26_GB00;
wire R10C37_X08;
wire R25C46_GBO0;
wire R12C36_GB00;
wire R15C37_GBO0;
wire R10C34_N82;
wire R28C46_D7;
wire R29C28_D6;
wire R28C19_W23;
wire R11C20_GB30;
wire R22C42_GB00;
wire R14C6_GT00;
wire R10C19_X05;
wire R18C17_GB10;
wire R4C9_GB40;
wire R26C30_GB50;
wire R22C34_GB50;
wire R27C42_GB30;
wire R8C36_GB10;
wire R9C19_GT00;
wire R14C42_GB30;
wire R10C43_Q4;
wire R27C23_GB20;
wire R21C1_GBO0;
wire R24C12_GT00;
wire R12C11_GBO1;
wire R7C32_GB20;
wire R23C42_GB70;
wire R4C4_GB00;
wire R10C25_C5;
wire R10C31_N81;
wire R6C40_GBO0;
wire R28C31_Q4;
wire R3C41_GB40;
wire R26C20_GB20;
wire R20C22_GBO1;
wire R1C28_Q3;
wire R28C46_W25;
wire R6C30_GT10;
wire R2C24_GB10;
wire R10C37_S83;
wire R16C13_GB00;
wire R10C27_C7;
wire R20C3_GB30;
wire R24C20_GB60;
wire R10C31_D4;
wire R3C3_GT10;
wire R26C14_GB60;
wire R3C3_GB40;
wire R14C9_GBO1;
wire R23C10_GT00;
wire R17C20_GBO1;
wire R20C40_SPINE24;
wire R28C22_LSR1;
wire R11C6_GB20;
wire R28C16_C2;
wire R4C27_GB70;
wire R17C6_GB20;
wire R21C19_GB40;
wire R20C33_GB50;
wire R10C19_W26;
wire R9C37_GB40;
wire R4C7_GT10;
wire R28C22_F4;
wire R22C25_GB60;
wire R8C12_GB00;
wire R23C19_GB10;
wire R10C37_X05;
wire R3C43_GB00;
wire R8C31_GT00;
wire R15C36_GBO1;
wire R13C35_GB60;
wire R20C26_SPINE18;
wire R17C5_GBO1;
wire R16C2_GB30;
wire R1C32_B4;
wire R10C13_X02;
wire R18C38_GB00;
wire R10C16_C1;
wire R23C30_GB30;
wire R2C2_GT10;
wire R3C14_GB70;
wire R9C2_GB60;
wire R18C22_GB60;
wire R28C31_W80;
wire R1C32_A1;
wire R24C30_GB40;
wire R5C25_GB70;
wire R21C30_GB20;
wire R10C28_E13;
wire R22C33_GB50;
wire R5C14_GT10;
wire R6C7_GB30;
wire R14C22_GB10;
wire R28C22_W12;
wire R6C14_GB20;
wire R15C10_GB30;
wire R15C45_GB10;
wire R10C19_A4;
wire R13C37_GB30;
wire R10C29_CE0;
wire R13C6_GT10;
wire R7C42_GB20;
wire R12C12_GB50;
wire R6C18_GB00;
wire R21C21_GB60;
wire R15C2_GB70;
wire R10C13_S82;
wire R18C20_GT00;
wire R10C22_E22;
wire R25C24_GB20;
wire R5C10_GBO1;
wire R21C42_GB70;
wire R28C43_Q7;
wire R24C31_GT00;
wire R22C18_GB00;
wire R10C28_F4;
wire R23C45_GB00;
wire R2C22_GBO1;
wire R7C23_GB60;
wire R26C24_GBO1;
wire R25C10_GB40;
wire R12C31_GT00;
wire R5C27_GB60;
wire R10C40_C4;
wire R24C25_GB70;
wire R10C16_E83;
wire R14C40_GT10;
wire R22C23_GB70;
wire R5C23_GB20;
wire R10C43_B4;
wire R20C24_GBO0;
wire R7C29_GB70;
wire R26C13_GB40;
wire R8C30_GBO0;
wire R5C14_GBO1;
wire R10C7_N26;
wire R14C21_GT00;
wire R10C22_X04;
wire R24C29_GB50;
wire R7C45_GB10;
wire R28C16_W11;
wire R28C4_C6;
wire R28C13_F2;
wire R13C24_GB40;
wire R9C26_GBO1;
wire R28C25_S10;
wire R6C42_GT10;
wire R1C1_X03;
wire R1C32_W27;
wire R25C25_GB50;
wire R11C23_GB10;
wire R6C15_GT00;
wire R26C16_GBO1;
wire R14C20_GB70;
wire R7C5_GB50;
wire R27C31_GB60;
wire R25C26_GT00;
wire R1C32_Q2;
wire R28C19_W12;
wire R3C29_GT00;
wire R5C37_GB40;
wire R18C32_GB70;
wire R10C26_E13;
wire R28C25_W26;
wire R26C32_GB30;
wire R1C47_B3;
wire R26C33_GB40;
wire R15C21_GB50;
wire R22C36_GB10;
wire R2C5_SPINE11;
wire R24C7_GB50;
wire R16C20_GB70;
wire R10C28_SPINE16;
wire R7C28_GB60;
wire R28C7_X07;
wire R23C20_GB30;
wire R21C11_GBO1;
wire R10C31_C0;
wire R13C12_GB50;
wire R26C42_GB30;
wire R10C16_S21;
wire R7C1_GT10;
wire R18C6_GBO1;
wire R28C28_EW10;
wire R10C43_W24;
wire R17C28_GB30;
wire R9C8_GBO1;
wire R9C11_GB50;
wire R10C43_E26;
wire R6C15_GB60;
wire R9C17_GB30;
wire R11C43_GB10;
wire R11C42_GT00;
wire R8C17_GB10;
wire R4C5_GT00;
wire R11C32_GB60;
wire R20C11_GB60;
wire R21C39_GB70;
wire R16C24_GB70;
wire R10C16_E82;
wire R11C15_GT10;
wire R10C19_C1;
wire R25C3_GB10;
wire R10C22_CE2;
wire R10C27_X05;
wire R8C30_GB30;
wire R10C28_C5;
wire R10C19_A5;
wire R28C34_SEL6;
wire R2C4_SPINE8;
wire R6C31_GB60;
wire R20C28_GT00;
wire R21C36_GB40;
wire R16C34_GB50;
wire R28C40_S83;
wire R14C44_GB70;
wire R10C34_Q6;
wire R18C26_GB10;
wire R24C27_GB30;
wire R11C25_GB50;
wire R15C39_GB00;
wire R27C33_GB50;
wire R10C10_C4;
wire R28C43_N25;
wire R2C34_GT00;
wire R3C15_GB70;
wire R20C31_GB50;
wire R6C30_GB50;
wire R4C38_GB00;
wire R10C27_UNK123;
wire R10C27_S26;
wire R10C28_E26;
wire R17C23_GB10;
wire R26C16_GB00;
wire R10C30_B2;
wire R17C32_GB10;
wire R27C34_GB70;
wire R20C36_GB40;
wire R10C37_E83;
wire R9C31_GB70;
wire R10C31_D3;
wire R8C7_GB00;
wire R16C43_GB20;
wire R28C22_B4;
wire R2C35_GB50;
wire R28C31_SN10;
wire R17C35_GB30;
wire R22C17_GB40;
wire R26C14_GB10;
wire R7C25_GT10;
wire R28C31_A5;
wire R10C22_S80;
wire R28C4_D1;
wire R10C30_W11;
wire R6C45_GB20;
wire R11C44_GB50;
wire R12C43_GBO0;
wire R8C6_GB40;
wire R4C25_GT00;
wire R28C46_N21;
wire R6C38_GB40;
wire R24C13_GBO1;
wire R10C37_E12;
wire R11C39_GB10;
wire R24C30_GT00;
wire R4C31_GB20;
wire R14C14_GB20;
wire R3C23_GBO1;
wire R15C33_GB60;
wire R20C28_GB20;
wire R10C16_E12;
wire R4C29_GB70;
wire R4C45_GB70;
wire R10C34_A2;
wire R10C29_SPINE24;
wire R21C18_GB10;
wire R2C6_GB00;
wire R11C45_GB50;
wire R28C40_F3;
wire R13C9_GB40;
wire R24C7_GB10;
wire R20C23_GBO0;
wire R16C41_GB00;
wire R10C19_EW10;
wire R28C43_C2;
wire R28C16_C5;
wire R10C16_C2;
wire R16C14_GBO0;
wire R13C36_GB40;
wire R4C22_GB20;
wire R16C17_GB00;
wire R28C19_X03;
wire R3C12_GBO0;
wire R18C11_GB40;
wire R10C29_A0;
wire R22C16_GT00;
wire R6C43_GBO1;
wire R18C46_GB00;
wire R1C47_SN10;
wire R28C28_E10;
wire R26C41_GBO0;
wire R15C10_GB00;
wire R2C13_GB20;
wire R14C10_GBO1;
wire R28C4_CLK2;
wire R26C27_GB00;
wire R3C34_GB00;
wire R6C34_GT10;
wire R8C39_GB40;
wire R6C29_GB00;
wire R3C33_GB60;
wire R9C43_GBO0;
wire R22C36_GB40;
wire R7C2_GB70;
wire R13C39_GBO0;
wire R10C31_CE1;
wire R5C21_GT10;
wire R6C22_GT00;
wire R6C35_GB40;
wire R10C19_S80;
wire R22C14_GB40;
wire R28C43_S26;
wire R2C16_GB20;
wire R11C27_GB00;
wire R3C43_GBO0;
wire R10C13_W11;
wire R25C42_GB70;
wire R27C11_GB60;
wire R3C30_GT10;
wire R10C26_F7;
wire R8C16_GB70;
wire R23C38_GBO0;
wire R17C4_GBO1;
wire R14C18_GB70;
wire R27C9_GBO1;
wire R22C31_GT00;
wire R22C44_GB60;
wire R24C13_GBO0;
wire R6C35_GT00;
wire R15C43_GT10;
wire R23C15_GBO0;
wire R15C13_GB00;
wire R15C25_GB70;
wire R3C3_GB60;
wire R10C28_S10;
wire R5C8_GT00;
wire R13C26_GB60;
wire R28C25_D3;
wire R2C12_SPINE8;
wire R9C37_GT00;
wire R3C45_GB30;
wire R17C22_GB20;
wire R15C38_GB20;
wire R12C39_GB50;
wire R28C34_Q4;
wire R29C28_E20;
wire R16C8_GT10;
wire R8C31_GB00;
wire R8C15_GB20;
wire R10C43_S82;
wire R29C28_A4;
wire R16C16_GB10;
wire R7C12_GB20;
wire R23C27_GB10;
wire R28C28_F6;
wire R28C19_E21;
wire R28C19_E13;
wire R20C22_GT00;
wire R17C20_GB10;
wire R7C26_GB20;
wire R10C37_S13;
wire R28C25_F0;
wire R24C25_GBO0;
wire R26C32_GBO1;
wire R25C15_GB20;
wire R23C15_GB30;
wire R13C10_GT10;
wire R27C42_GT00;
wire R3C24_GB40;
wire R22C14_GB60;
wire R10C31_Q7;
wire R10C37_SEL2;
wire R1C28_N25;
wire R28C4_C1;
wire R11C3_GBO1;
wire R28C10_SEL7;
wire R28C46_SN20;
wire R15C8_GBO1;
wire R10C30_SPINE0;
wire R5C16_GB50;
wire R28C28_F0;
wire R20C44_GB60;
wire R20C42_GB20;
wire R1C32_Q5;
wire R28C31_B3;
wire R8C44_GB30;
wire R28C25_N81;
wire R2C18_GBO1;
wire R20C10_GB00;
wire R9C34_GBO0;
wire R10C40_B0;
wire R28C40_N27;
wire R20C22_GB60;
wire R27C29_GT10;
wire R15C29_GB00;
wire R27C17_GT10;
wire R10C19_W10;
wire R10C40_E11;
wire R14C16_GB70;
wire R11C12_GT00;
wire R16C25_GB30;
wire R25C7_GBO1;
wire R22C23_GB60;
wire R16C18_GB10;
wire R15C19_GB40;
wire R6C4_GB40;
wire R6C8_GB60;
wire R15C13_GT10;
wire R14C16_GB10;
wire R15C12_GB50;
wire R13C3_GB50;
wire R13C5_GBO1;
wire R28C37_S20;
wire R8C25_GB30;
wire R13C23_GBO0;
wire R10C27_B6;
wire R22C34_GB40;
wire R6C26_GB60;
wire R18C35_GB20;
wire R28C7_E80;
wire R11C24_GBO0;
wire R11C3_GB50;
wire R1C47_F7;
wire R2C6_GB10;
wire R22C3_GB40;
wire R25C10_GB60;
wire R21C22_GB70;
wire R1C32_F5;
wire R11C24_GT00;
wire R28C22_S11;
wire R9C43_GB70;
wire R2C13_GB70;
wire R28C31_S20;
wire R7C19_GB50;
wire R18C37_GT10;
wire R10C37_SEL0;
wire R9C6_GB10;
wire R24C15_GB10;
wire R22C2_GBO1;
wire R20C40_GT00;
wire R9C37_GB70;
wire R8C2_GB10;
wire R10C27_Q4;
wire R15C38_GB50;
wire R10C27_D1;
wire R8C27_GBO1;
wire R14C16_GT00;
wire R24C38_GB50;
wire R3C11_GT00;
wire R25C38_GB40;
wire R11C41_GB40;
wire R22C23_GBO1;
wire R8C41_GB70;
wire R11C7_GB00;
wire R6C32_GB10;
wire R16C32_GB10;
wire R28C31_D1;
wire R6C30_GB20;
wire R14C19_GB60;
wire R12C11_GB70;
wire R15C24_GBO0;
wire R17C2_GB50;
wire R6C31_GBO0;
wire R6C45_GB30;
wire R10C43_E23;
wire R18C22_GB00;
wire R27C36_GT00;
wire R28C16_D5;
wire R9C2_GB00;
wire R24C4_GT10;
wire R10C28_N12;
wire R10C16_X01;
wire R27C18_GT00;
wire R4C38_GT00;
wire R23C7_GB00;
wire R18C43_GB70;
wire R28C10_E13;
wire R11C26_GBO0;
wire R10C22_C5;
wire R29C28_SEL7;
wire R28C25_N21;
wire R20C5_GB40;
wire R28C37_CE2;
wire R5C18_GB00;
wire R28C31_E12;
wire R26C11_GB70;
wire R21C40_GB40;
wire R22C14_GB30;
wire R28C40_S26;
wire R26C43_GB20;
wire R13C19_GBO0;
wire R6C36_GB30;
wire R15C45_GBO1;
wire R17C34_GB30;
wire R10C37_SEL7;
wire R28C34_SEL1;
wire R7C31_GBO1;
wire R28C34_N20;
wire R6C6_GB70;
wire R3C4_GT00;
wire R16C16_GB30;
wire R10C40_SEL5;
wire R6C4_GB70;
wire R9C22_GB30;
wire R22C21_GBO0;
wire R1C47_B1;
wire R10C27_E24;
wire R28C28_E13;
wire R10C31_C3;
wire R12C27_GT00;
wire R18C36_GT10;
wire R11C20_GBO1;
wire R4C29_GB00;
wire R16C37_GB60;
wire R10C26_E80;
wire R5C32_GT10;
wire R24C2_GBO1;
wire R12C9_GB70;
wire R16C45_GB70;
wire R5C9_GT10;
wire R28C19_X04;
wire R23C6_GT10;
wire R20C30_GBO0;
wire R18C41_GB30;
wire R26C8_GB30;
wire R17C12_GB60;
wire R2C45_GB70;
wire R5C20_GT00;
wire R23C19_GB30;
wire R25C36_GBO1;
wire R1C28_E24;
wire R8C8_GB00;
wire R28C4_D7;
wire R12C27_GB10;
wire R25C37_GB70;
wire R28C25_S82;
wire R9C33_GB50;
wire R10C40_E27;
wire R24C9_GB40;
wire R7C24_GT00;
wire R9C5_GB70;
wire R17C24_GB70;
wire R8C39_GB20;
wire R26C44_GB30;
wire R23C37_GB60;
wire R21C12_GB70;
wire R22C8_GB50;
wire R14C43_GB40;
wire R25C9_GB00;
wire R15C4_GB40;
wire R10C7_W82;
wire R17C6_GBO0;
wire R6C29_GBO0;
wire R18C8_GT00;
wire R8C14_GB60;
wire R17C39_GB40;
wire R10C13_A7;
wire R10C19_SN20;
wire R26C26_GT00;
wire R10C28_LSR1;
wire R17C25_GT10;
wire R28C4_N24;
wire R2C12_GT10;
wire R4C19_GB00;
wire R5C4_GB60;
wire R22C4_GBO0;
wire R13C41_GT00;
wire R6C31_GT00;
wire R10C10_S21;
wire R10C16_EW20;
wire R25C32_GB40;
wire R11C27_GT00;
wire R17C36_GB20;
wire R10C26_D1;
wire R10C37_A4;
wire R4C14_GT10;
wire R8C26_GB00;
wire R28C46_W26;
wire R8C9_GB10;
wire R28C37_E23;
wire R20C30_GB70;
wire R7C13_GB10;
wire R29C28_N24;
wire R11C3_GB30;
wire R24C42_GB20;
wire R6C37_GB30;
wire R10C7_D6;
wire R28C37_EW10;
wire R13C36_GT10;
wire R21C40_GT10;
wire R10C37_A3;
wire R26C4_GT00;
wire R6C25_GB70;
wire R12C8_GT10;
wire R2C42_GT10;
wire R12C35_GT00;
wire R21C14_GB50;
wire R9C45_GB50;
wire R17C41_GB40;
wire R27C42_GBO1;
wire R23C18_GB60;
wire R15C16_GT00;
wire R24C35_GB70;
wire R3C2_GT00;
wire R9C28_GB20;
wire R10C30_SEL1;
wire R16C8_GB20;
wire R28C31_D2;
wire R12C14_GB00;
wire R13C39_GT10;
wire R28C37_B5;
wire R3C42_GB70;
wire R3C8_GB30;
wire R14C17_GB70;
wire R10C30_CLK0;
wire R28C16_F5;
wire R16C4_GB30;
wire R27C37_GT00;
wire R18C19_GB60;
wire R14C23_GT00;
wire R2C7_GB30;
wire R21C28_GT00;
wire R7C36_GB00;
wire R22C38_GB10;
wire R25C34_GB40;
wire R4C41_GB70;
wire R15C2_GB60;
wire R1C1_A2;
wire R10C40_A1;
wire R29C28_SN10;
wire R17C11_GB20;
wire R17C9_GBO1;
wire R26C2_GBO1;
wire R2C10_GT10;
wire R1C47_SEL6;
wire R5C15_GB70;
wire R10C40_CLK1;
wire R21C38_GB30;
wire R28C7_N10;
wire R20C9_GBO0;
wire R28C25_E21;
wire R6C18_GB30;
wire R18C14_GT00;
wire R12C2_GB00;
wire R10C30_SEL4;
wire R10C43_F0;
wire R14C26_GT10;
wire R11C23_GB70;
wire R7C33_GB70;
wire R9C39_GB70;
wire R28C28_N81;
wire R10C34_LSR0;
wire R24C46_GT00;
wire R10C10_SEL1;
wire R10C10_D2;
wire R2C18_GT00;
wire R9C38_GBO1;
wire R2C5_GB10;
wire R8C24_GB20;
wire R28C16_N10;
wire R26C40_GB10;
wire R12C18_GB60;
wire R28C28_CE0;
wire R18C29_GBO1;
wire R8C24_GBO1;
wire R10C22_SEL6;
wire R21C38_GT10;
wire R8C20_GBO1;
wire R10C31_A2;
wire R9C44_GB70;
wire R12C4_GB00;
wire R12C23_GB30;
wire R11C21_GB40;
wire R1C1_CLK0;
wire R16C29_GT00;
wire R1C28_N80;
wire R12C9_GB30;
wire R9C35_GB70;
wire R28C34_X04;
wire R4C4_GB70;
wire R7C35_GB60;
wire R24C16_GBO0;
wire R1C1_D3;
wire R11C3_GB60;
wire R4C39_GB70;
wire R20C17_GT00;
wire R18C19_GB70;
wire R13C10_GB50;
wire R25C38_GT10;
wire R1C32_A0;
wire R22C8_GB00;
wire R28C37_A5;
wire R7C26_GB70;
wire R18C43_GB30;
wire R1C1_S21;
wire R15C30_GB20;
wire R3C16_GT00;
wire R18C25_GB50;
wire R6C16_GT10;
wire R27C3_GT00;
wire R1C28_D6;
wire R26C12_GB40;
wire R27C24_GT00;
wire R28C31_E24;
wire R21C8_GBO0;
wire R11C8_GB00;
wire R18C32_GB00;
wire R28C40_N13;
wire R25C25_GB10;
wire R20C42_GB60;
wire R10C13_S80;
wire R23C38_GBO1;
wire R23C19_GB00;
wire R1C28_C2;
wire R21C35_GT00;
wire R28C19_S20;
wire R9C15_GT10;
wire R4C7_GB60;
wire R28C46_W82;
wire R20C45_GB10;
wire R14C45_GB40;
wire R22C20_GB20;
wire R14C36_GT00;
wire R6C27_GT00;
wire R3C14_GB40;
wire R24C2_GB70;
wire R11C40_GB60;
wire R28C40_S23;
wire R10C25_N11;
wire R10C27_D0;
wire R24C19_GB00;
wire R3C8_GT10;
wire R14C16_GT10;
wire R20C35_GB00;
wire R8C6_GB00;
wire R17C31_GB40;
wire R17C27_GBO1;
wire R11C14_GB20;
wire R20C42_GT10;
wire R10C27_LSR1;
wire R8C41_GBO0;
wire R26C17_GT10;
wire R24C4_GBO0;
wire R24C2_GB50;
wire R14C29_GB10;
wire R14C3_GT10;
wire R17C20_GB00;
wire R22C45_GB40;
wire R28C25_SN20;
wire R20C32_GB60;
wire R28C43_A2;
wire R24C37_GB50;
wire R28C10_S80;
wire R12C42_GB30;
wire R20C13_SPINE19;
wire R10C31_Q4;
wire R6C30_GB40;
wire R10C22_B5;
wire R24C4_GB30;
wire R26C21_GB40;
wire R6C2_GB20;
wire R8C3_GB00;
wire R14C10_GB00;
wire R13C26_GB30;
wire R20C35_GB30;
wire R26C15_GB00;
wire R22C25_GB30;
wire R13C41_GB50;
wire R25C26_GB20;
wire R10C40_E23;
wire R28C40_E25;
wire R28C40_S12;
wire R1C47_E20;
wire R10C13_S23;
wire R18C11_GB00;
wire R7C30_GB50;
wire R27C45_GB60;
wire R25C45_GT10;
wire R5C39_GB10;
wire R29C28_W13;
wire R23C9_GB10;
wire R10C26_B5;
wire R13C11_GB50;
wire R5C8_GB40;
wire R16C15_GT00;
wire R20C4_GT00;
wire R13C18_GBO0;
wire R4C38_GB20;
wire R14C33_GBO1;
wire R5C3_GB00;
wire R7C33_GB00;
wire R10C30_S83;
wire R1C28_E26;
wire R5C21_GT00;
wire R16C14_GBO1;
wire R28C13_B0;
wire R28C16_D6;
wire R6C4_GB50;
wire R14C25_GT00;
wire R20C3_GB40;
wire R6C43_GB50;
wire R15C40_GT10;
wire R10C30_X03;
wire R15C22_GBO0;
wire R18C37_GBO0;
wire R12C8_GB10;
wire R27C17_GB70;
wire R7C17_GT00;
wire R14C33_GB30;
wire R24C43_GB00;
wire R22C22_GB60;
wire R1C47_Q0;
wire R12C46_GBO1;
wire R14C26_GB00;
wire R10C29_E83;
wire R28C10_F0;
wire R6C37_GB00;
wire R5C45_GT10;
wire R4C5_GB20;
wire R6C16_GB60;
wire R2C41_GB30;
wire R21C33_GB70;
wire R28C31_A4;
wire R28C46_B7;
wire R12C35_GB30;
wire R1C47_CLK1;
wire R22C24_GB20;
wire R28C10_B1;
wire R16C46_GBO0;
wire R11C8_GB50;
wire R17C37_GB10;
wire R28C28_SN20;
wire R6C36_GB40;
wire R11C25_GBO0;
wire R28C31_Q7;
wire R28C31_N10;
wire R10C30_D5;
wire R8C43_GB10;
wire R16C34_GB60;
wire R21C9_GB60;
wire R14C16_GBO1;
wire R28C46_CE1;
wire R3C4_GB00;
wire R20C13_GT10;
wire R2C15_GB10;
wire R25C44_GT00;
wire R22C35_GB70;
wire R10C25_Q5;
wire R29C28_EW20;
wire R7C9_GT00;
wire R2C28_GB20;
wire R22C44_GB70;
wire R10C43_N13;
wire R13C18_GB20;
wire R27C11_GB10;
wire R15C41_GBO0;
wire R15C3_GB00;
wire R27C11_GB50;
wire R11C32_GB30;
wire R17C9_GBO0;
wire R15C2_GBO0;
wire R10C19_SEL6;
wire R28C22_B7;
wire R14C12_GB30;
wire R11C6_GB40;
wire R20C27_GBO1;
wire R10C25_N27;
wire R6C43_GB70;
wire R10C29_D6;
wire R16C40_GT00;
wire R10C22_N27;
wire R21C24_GB50;
wire R5C13_GT10;
wire R10C7_N10;
wire R10C26_W13;
wire R10C37_X02;
wire R28C13_A5;
wire R10C30_UNK123;
wire R4C6_GB50;
wire R8C19_GB60;
wire R27C10_GB00;
wire R28C37_C1;
wire R23C29_GT00;
wire R1C47_C4;
wire R25C18_GT10;
wire R18C7_GB70;
wire R27C10_GT00;
wire R12C6_GB00;
wire R13C40_GB50;
wire R23C36_GB60;
wire R25C14_GBO0;
wire R10C16_D1;
wire R2C38_GBO0;
wire R28C10_B5;
wire R20C38_GBO0;
wire R5C2_GT10;
wire R4C11_GT10;
wire R13C45_GB60;
wire R10C26_N27;
wire R14C21_GBO1;
wire R28C46_B0;
wire R20C24_GT00;
wire R1C32_X02;
wire R14C44_GBO1;
wire R15C3_GB50;
wire R10C43_N21;
wire R28C34_LSR2;
wire R20C4_GB60;
wire R9C18_GB30;
wire R7C44_GBO1;
wire R4C34_GB70;
wire R16C9_GBO1;
wire R22C3_GBO0;
wire R8C21_GB70;
wire R28C34_E10;
wire R10C43_S20;
wire R13C8_GB60;
wire R17C38_GB50;
wire R18C16_GB20;
wire R21C10_GBO0;
wire R13C23_GB40;
wire R10C19_D1;
wire R27C15_GT10;
wire R27C40_GB10;
wire R28C10_E80;
wire R22C39_GT00;
wire R17C5_GB00;
wire R12C22_GB10;
wire R24C3_GT00;
wire R12C30_GB40;
wire R12C19_GBO0;
wire R6C42_GB40;
wire R21C35_GBO1;
wire R10C10_E22;
wire R10C26_X08;
wire R15C44_GB40;
wire R28C34_F1;
wire R22C14_GB70;
wire R3C24_GBO1;
wire R10C13_N21;
wire R29C28_N20;
wire R5C45_GB00;
wire R10C25_E26;
wire R17C42_GB50;
wire R26C32_GB20;
wire R1C28_W20;
wire R10C26_W10;
wire R10C37_SEL6;
wire R15C38_GT10;
wire R3C10_GB70;
wire R14C31_GBO0;
wire R10C26_D3;
wire R27C25_GB60;
wire R12C14_GB50;
wire R15C12_GT10;
wire R12C10_GB10;
wire R14C21_GT10;
wire R28C40_W10;
wire R26C24_GB60;
wire R24C46_GB20;
wire R5C45_GB20;
wire R10C25_N12;
wire R10C16_C7;
wire R28C4_D3;
wire R23C26_GB60;
wire R13C27_GB70;
wire R18C34_GB60;
wire R1C47_A6;
wire R28C10_E25;
wire R10C10_SEL6;
wire R26C44_GT10;
wire R15C21_GB10;
wire R13C5_GB00;
wire R4C40_GT10;
wire R6C44_GT00;
wire R10C25_X01;
wire R10C29_W13;
wire R28C22_SEL0;
wire R3C31_GB30;
wire R28C34_B1;
wire R15C21_GT10;
wire R29C28_X06;
wire R14C26_GBO0;
wire R9C12_GT00;
wire R11C39_GB00;
wire R11C46_GB10;
wire R7C32_GT10;
wire R3C44_GB40;
wire R6C25_GBO1;
wire R8C24_GB30;
wire R15C12_GB20;
wire R10C10_N22;
wire R21C4_GT00;
wire R3C24_GBO0;
wire R28C22_W11;
wire R28C19_Q2;
wire R25C28_GB20;
wire R16C10_GBO1;
wire R28C37_D0;
wire R14C20_GT10;
wire R20C11_GB10;
wire R25C19_GB30;
wire R15C32_GBO1;
wire R28C19_E11;
wire R20C37_GT00;
wire R21C27_GBO1;
wire R10C10_A6;
wire R1C28_W12;
wire R16C43_GB00;
wire R23C7_GBO0;
wire R21C3_GB60;
wire R4C35_GB50;
wire R28C37_C5;
wire R28C10_LSR0;
wire R10C29_E20;
wire R23C23_GT00;
wire R8C6_GBO0;
wire R9C28_GT00;
wire R16C11_GB60;
wire R5C31_GBO0;
wire R10C22_CLK1;
wire R21C38_GBO0;
wire R22C42_GB10;
wire R28C40_N26;
wire R3C19_GT00;
wire R28C7_S13;
wire R13C14_GBO0;
wire R25C28_GB50;
wire R24C35_GB30;
wire R2C22_SPINE10;
wire R12C25_GB60;
wire R27C44_GB70;
wire R10C7_LSR1;
wire R28C4_C0;
wire R28C31_W82;
wire R26C30_GB30;
wire R9C24_GB30;
wire R13C42_GB40;
wire R4C30_GT10;
wire R20C3_GT00;
wire R4C26_GB40;
wire R1C1_B0;
wire R4C29_GB10;
wire R28C16_A6;
wire R28C28_SN10;
wire R14C27_GB40;
wire R14C5_GB10;
wire R24C27_GB40;
wire R9C1_GBO0;
wire R10C10_W80;
wire R10C29_D3;
wire R3C14_GB60;
wire R28C13_W21;
wire R28C34_W22;
wire R15C18_GB20;
wire R20C7_SPINE21;
wire R12C22_GB60;
wire R5C22_GB60;
wire R6C22_GB70;
wire R17C43_GBO0;
wire R28C4_D5;
wire R28C25_W13;
wire R3C46_GT00;
wire R20C37_GBO0;
wire R10C22_W83;
wire R25C8_GBO1;
wire R7C10_GT00;
wire R24C5_GB40;
wire R6C42_GB30;
wire R10C26_S25;
wire R13C11_GB30;
wire R28C43_N20;
wire R1C47_W12;
wire R13C23_GB50;
wire R10C13_W26;
wire R10C43_CLK1;
wire R21C11_GB20;
wire R7C43_GB30;
wire R5C23_GB70;
wire R28C43_S81;
wire R28C19_B3;
wire R6C43_GB60;
wire R14C22_GB00;
wire R2C24_SPINE8;
wire R8C7_GBO1;
wire R10C7_E20;
wire R10C29_LSR1;
wire R28C10_E27;
wire R26C9_GBO1;
wire R8C31_GB30;
wire R28C28_W82;
wire R29C28_D0;
wire R28C22_SEL3;
wire R10C26_X03;
wire R24C36_GB40;
wire R28C19_B4;
wire R13C40_GB20;
wire R21C14_GBO1;
wire R21C21_GT10;
wire R18C6_GB30;
wire R11C41_GT10;
wire R1C1_E12;
wire R29C28_D5;
wire R20C23_GB30;
wire R3C24_GT10;
wire R10C10_E10;
wire R28C28_E81;
wire R28C25_S25;
wire R10C13_W20;
wire R14C38_GT10;
wire R22C41_GT10;
wire R28C28_S26;
wire R20C12_GB20;
wire R24C24_GB00;
wire R10C25_F6;
wire R6C25_GBO0;
wire R8C26_GB60;
wire R25C23_GB20;
wire R28C40_C1;
wire R27C8_GB10;
wire R10C34_A1;
wire R1C1_C2;
wire R1C1_CE0;
wire R13C10_GB10;
wire R28C10_E81;
wire R4C32_GB00;
wire R2C14_GT10;
wire R16C24_GB30;
wire R10C43_C2;
wire R14C21_GB70;
wire R23C4_GB70;
wire R28C7_B7;
wire R13C26_GB50;
wire R14C33_GB20;
wire R5C13_GB00;
wire R21C30_GB60;
wire R1C32_X03;
wire R7C33_GB30;
wire R14C23_GB40;
wire R9C7_GBO0;
wire R17C10_GB00;
wire R18C29_GB60;
wire R26C23_GBO0;
wire R3C16_GBO0;
wire R12C11_GB30;
wire R4C15_GB50;
wire R27C33_GB00;
wire R22C37_GB00;
wire R28C13_S21;
wire R28C37_Q4;
wire R7C4_GT10;
wire R1C28_X08;
wire R8C2_GB30;
wire R18C21_GB40;
wire R16C22_GB60;
wire R17C43_GT10;
wire R3C42_GB40;
wire R20C39_GB30;
wire R20C44_SPINE24;
wire R14C9_GB20;
wire R27C1_GT00;
wire R22C46_GB50;
wire R5C25_GT10;
wire R5C18_GB40;
wire R6C34_GB60;
wire R8C39_GT00;
wire R4C43_GB30;
wire R14C32_GBO0;
wire R28C13_W22;
wire R6C31_GB40;
wire R12C4_GBO0;
wire R28C43_S20;
wire R13C6_GB70;
wire R12C37_GB00;
wire R26C13_GBO1;
wire R8C27_GB60;
wire R18C42_GB00;
wire R18C29_GB00;
wire R28C46_X08;
wire R1C28_N83;
wire R10C13_B1;
wire R12C15_GBO1;
wire R18C38_GT10;
wire R27C21_GT00;
wire R13C23_GB10;
wire R13C41_GB00;
wire R4C16_GB70;
wire R26C42_GB50;
wire R3C12_GB30;
wire R10C43_D1;
wire R24C40_GBO1;
wire R10C22_D4;
wire R28C4_Q7;
wire R14C12_GBO1;
wire R13C16_GB10;
wire R28C25_E22;
wire R14C15_GB00;
wire R14C29_GB50;
wire R8C28_GB60;
wire R9C46_GBO0;
wire R10C10_C6;
wire R28C16_B3;
wire R8C5_GB00;
wire R22C27_GBO0;
wire R10C29_B7;
wire R9C11_GB70;
wire R17C6_GB10;
wire R25C36_GT00;
wire R7C24_GB40;
wire R16C29_GB40;
wire R18C41_GBO1;
wire R22C19_GBO0;
wire R28C7_S12;
wire R20C3_GB20;
wire R23C17_GBO1;
wire R2C11_GBO1;
wire R4C9_GB30;
wire R10C27_D2;
wire R1C47_S82;
wire R12C38_GT10;
wire R2C41_GB00;
wire R26C40_GB00;
wire R10C40_X07;
wire R28C4_W83;
wire R16C45_GT00;
wire R28C46_W81;
wire R7C15_GB60;
wire R28C4_Q1;
wire R10C37_SEL5;
wire R5C9_GB10;
wire R10C27_S22;
wire R13C29_GB60;
wire R17C3_GT10;
wire R22C23_GT00;
wire R28C37_S24;
wire R4C25_GT10;
wire R15C36_GT00;
wire R16C45_GT10;
wire R11C36_GB30;
wire R3C23_GB70;
wire R25C42_GB20;
wire R18C37_GB40;
wire R2C27_GB60;
wire R25C31_GB50;
wire R10C7_W27;
wire R3C18_GB20;
wire R28C13_B7;
wire R28C25_F5;
wire R28C31_S82;
wire R3C39_GB20;
wire R11C5_GB10;
wire R9C21_GBO1;
wire R20C6_GBO1;
wire R1C32_Q1;
wire R5C38_GT10;
wire R3C42_GB10;
wire R27C7_GB30;
wire R10C25_A4;
wire R10C43_N27;
wire R16C20_GB00;
wire R4C42_GB10;
wire R10C10_B2;
wire R10C43_X01;
wire R14C6_GB00;
wire R2C32_GB10;
wire R24C37_GB30;
wire R28C22_E25;
wire R23C8_GT10;
wire R10C19_CLK1;
wire R9C35_GB10;
wire R13C35_GT00;
wire R17C17_GB10;
wire R28C22_D1;
wire R9C26_GBO0;
wire R12C40_GBO1;
wire R14C10_GB50;
wire R9C40_GB60;
wire R16C30_GB10;
wire R29C28_A6;
wire R24C31_GBO0;
wire R3C6_GB50;
wire R3C3_GT00;
wire R27C37_GB60;
wire R25C26_GB40;
wire R21C9_GBO0;
wire R26C41_GT10;
wire R23C32_GT10;
wire R21C3_GB50;
wire R27C36_GB60;
wire R10C34_SEL2;
wire R10C31_D1;
wire R16C33_GBO0;
wire R28C37_E24;
wire R8C44_GB40;
wire R24C3_GB10;
wire R5C16_GB60;
wire R26C7_GBO0;
wire R14C9_GB50;
wire R21C19_GB00;
wire R27C25_GB50;
wire R18C3_GB70;
wire R8C44_GB60;
wire R28C4_C5;
wire R29C28_W12;
wire R28C43_X06;
wire R23C21_GB00;
wire R17C44_GB40;
wire R23C43_GT00;
wire R26C46_GB30;
wire R3C3_GB50;
wire R21C40_GBO1;
wire R20C23_GB20;
wire R4C6_GB10;
wire R14C46_GB70;
wire R10C29_N26;
wire R20C19_GB50;
wire R27C21_GB30;
wire R16C6_GBO0;
wire R27C18_GBO1;
wire R8C44_GB50;
wire R16C26_GB00;
wire R24C9_GBO0;
wire R10C27_N81;
wire R24C28_GB00;
wire R18C13_GB40;
wire R5C4_GT10;
wire R3C28_GB30;
wire R12C11_GT10;
wire R3C46_GB50;
wire R1C28_B1;
wire R28C34_X05;
wire R18C5_GT10;
wire R13C40_GB70;
wire R25C37_GB30;
wire R4C24_GT10;
wire R10C19_E81;
wire R10C25_D1;
wire R10C43_W21;
wire R4C15_GB10;
wire R23C25_GB20;
wire R24C22_GBO0;
wire R14C46_GB40;
wire R10C26_X01;
wire R1C32_A6;
wire R28C16_A7;
wire R9C26_GB00;
wire R27C42_GB10;
wire R12C38_GBO1;
wire R1C32_S22;
wire R10C30_N11;
wire R12C42_GT00;
wire R22C28_GB60;
wire R23C43_GT10;
wire R27C6_GB10;
wire R13C16_GB40;
wire R5C40_GT10;
wire R22C6_GB00;
wire R25C4_GB10;
wire R26C27_GT00;
wire R17C14_GB20;
wire R28C34_CE1;
wire R10C34_S23;
wire R10C10_W12;
wire R28C31_CLK0;
wire R23C6_GT00;
wire R7C19_GB40;
wire R10C40_W13;
wire R27C13_GB00;
wire R9C29_GB60;
wire R15C21_GB40;
wire R8C15_GT10;
wire R10C31_S13;
wire R9C3_GB40;
wire R25C4_GB50;
wire R4C34_GB40;
wire R6C8_GT00;
wire R22C3_GB00;
wire R28C40_W21;
wire R9C34_GB50;
wire R28C43_X02;
wire R18C12_GB40;
wire R14C30_GB30;
wire R23C21_GBO1;
wire R10C31_E22;
wire R28C34_W13;
wire R24C11_GBO0;
wire R17C8_GB30;
wire R5C45_GBO1;
wire R14C15_GBO0;
wire R28C19_C2;
wire R18C7_GB00;
wire R13C15_GT10;
wire R6C27_GBO1;
wire R16C12_GB20;
wire R13C19_GB20;
wire R25C20_GB70;
wire R1C28_C0;
wire R23C13_GB10;
wire R21C11_GB10;
wire R17C7_GBO1;
wire R14C28_GB60;
wire R10C29_SEL2;
wire R10C10_B1;
wire R2C8_GB60;
wire R15C17_GB30;
wire R9C7_GBO1;
wire R28C22_A6;
wire R10C43_SEL5;
wire R1C1_C1;
wire R5C16_GB20;
wire R28C4_F1;
wire R29C28_S82;
wire R10C22_D2;
wire R27C41_GB20;
wire R18C9_GB70;
wire R10C34_D6;
wire R9C33_GBO1;
wire R10C30_E21;
wire R22C2_GB20;
wire R24C22_GB50;
wire R6C25_GB30;
wire R27C22_GB10;
wire R22C32_GB20;
wire R17C1_GT00;
wire R10C43_E21;
wire R28C7_X01;
wire R13C28_GB10;
wire R22C38_GB00;
wire R18C39_GT00;
wire R17C25_GBO0;
wire R13C2_GB20;
wire R15C39_GB10;
wire R10C40_N12;
wire R13C21_GB40;
wire R28C19_W26;
wire R27C29_GB20;
wire R6C8_GB30;
wire R23C37_GBO0;
wire R10C26_B7;
wire R23C17_GT10;
wire R25C33_GB70;
wire R14C2_GBO1;
wire R17C11_GT00;
wire R8C42_GT10;
wire R9C30_GT10;
wire R20C13_GB10;
wire R23C9_GBO0;
wire R17C32_GB30;
wire R5C46_GBO0;
wire R1C28_B4;
wire R23C32_GB30;
wire R10C40_E83;
wire R13C15_GB00;
wire R28C7_W83;
wire R28C46_A5;
wire R10C22_SEL4;
wire R10C29_X04;
wire R17C4_GB70;
wire R3C13_GB30;
wire R25C21_GB30;
wire R1C32_F6;
wire R10C34_D1;
wire R28C37_B3;
wire R26C4_GB40;
wire R8C13_GT10;
wire R4C44_GB70;
wire R15C11_GB40;
wire R26C38_GB60;
wire R21C17_GB70;
wire R10C37_N25;
wire R11C11_GT10;
wire R20C20_GBO1;
wire R25C27_GB60;
wire R22C10_GB60;
wire R21C11_GB60;
wire R2C32_GT10;
wire R28C4_S23;
wire R13C36_GB60;
wire R17C21_GB10;
wire R17C16_GB00;
wire R10C37_D6;
wire R18C16_GB50;
wire R28C40_Q7;
wire R24C30_GBO0;
wire R10C34_CE1;
wire R18C36_GB50;
wire R6C46_GB30;
wire R6C2_GB60;
wire R28C16_B5;
wire R13C25_GT10;
wire R24C14_GT10;
wire R18C27_GBO1;
wire R4C32_GB50;
wire R15C41_GT00;
wire R21C7_GBO1;
wire R24C18_GT00;
wire R24C31_GB70;
wire R8C34_GT10;
wire R4C17_GB70;
wire R10C27_W12;
wire R20C12_SPINE20;
wire R1C1_E21;
wire R15C15_GB20;
wire R23C35_GB00;
wire R24C13_GB50;
wire R12C15_GB10;
wire R3C14_GT00;
wire R10C10_Q3;
wire R11C7_GB10;
wire R5C2_GB70;
wire R14C24_GB70;
wire R9C37_GB20;
wire R15C44_GB20;
wire R23C17_GB50;
wire R23C18_GB50;
wire R28C37_W12;
wire R18C20_GB10;
wire R10C19_E26;
wire R27C31_GB70;
wire R24C10_GB10;
wire R16C46_GT10;
wire R20C25_GB20;
wire R9C40_GB30;
wire R1C28_W81;
wire R10C7_E13;
wire R28C37_Q1;
wire R5C17_GT00;
wire R18C12_GT10;
wire R2C7_GB10;
wire R9C7_GB10;
wire R28C31_S13;
wire R8C33_GB10;
wire R17C13_GB50;
wire R18C37_GB50;
wire R1C1_W11;
wire R4C14_GT00;
wire R14C6_GT10;
wire R1C32_B6;
wire R11C30_GB10;
wire R25C32_GT00;
wire R29C28_C6;
wire R7C4_GBO0;
wire R10C13_E82;
wire R10C31_W22;
wire R23C10_GB70;
wire R2C46_GT10;
wire R7C1_GBO0;
wire R4C42_GB00;
wire R28C19_D4;
wire R28C46_F2;
wire R28C37_W24;
wire R28C13_SEL2;
wire R2C32_GT00;
wire R15C24_GB70;
wire R6C22_GB00;
wire R13C42_GBO1;
wire R10C30_N26;
wire R1C28_N20;
wire R28C13_Q5;
wire R28C28_S12;
wire R13C33_GB40;
wire R28C40_S25;
wire R6C13_GB50;
wire R11C12_GB30;
wire R23C15_GB40;
wire R10C29_E26;
wire R9C46_GB60;
wire R21C7_GB00;
wire R17C5_GBO0;
wire R28C34_N11;
wire R16C21_GB00;
wire R28C16_E83;
wire R2C18_SPINE10;
wire R24C33_GB10;
wire R8C37_GB60;
wire R24C32_GB30;
wire R26C45_GB40;
wire R29C28_E27;
wire R2C41_GT00;
wire R23C34_GB20;
wire R21C28_GT10;
wire R10C31_E12;
wire R5C32_GBO1;
wire R10C7_D0;
wire R1C47_S10;
wire R29C28_N25;
wire R4C19_GBO0;
wire R28C25_LSR0;
wire R15C7_GB70;
wire R10C28_E83;
wire R22C35_GT10;
wire R17C35_GB50;
wire R21C40_GB70;
wire R10C25_F4;
wire R5C25_GBO1;
wire R22C39_GT10;
wire R26C34_GB00;
wire R20C14_GB40;
wire R24C2_GB40;
wire R12C29_GB30;
wire R25C40_GB30;
wire R22C8_GT10;
wire R18C6_GT10;
wire R22C11_GB40;
wire R24C46_GB30;
wire R25C13_GBO1;
wire R28C7_W23;
wire R9C34_GB00;
wire R10C16_S11;
wire R26C3_GT10;
wire R23C33_GB00;
wire R11C34_GB40;
wire R10C22_F5;
wire R25C9_GB50;
wire R16C7_GT00;
wire R23C19_GB60;
wire R17C40_GB30;
wire R28C31_X07;
wire R23C38_GB10;
wire R9C29_GBO1;
wire R1C1_SN10;
wire R20C36_GT10;
wire R28C37_N25;
wire R7C23_GB70;
wire R22C30_GB30;
wire R21C30_GT10;
wire R6C5_GB10;
wire R6C34_GB50;
wire R10C7_A0;
wire R2C19_GT00;
wire R10C10_Q6;
wire R10C10_D3;
wire R7C13_GB50;
wire R5C6_GB30;
wire R24C11_GB30;
wire R4C30_GB40;
wire R10C19_S10;
wire R28C10_SN20;
wire R22C17_GT10;
wire R22C3_GB20;
wire R6C25_GB50;
wire R16C7_GB70;
wire R13C34_GB00;
wire R10C13_S27;
wire R28C28_D2;
wire R28C4_N12;
wire R10C19_C7;
wire R10C25_X06;
wire R13C7_GB50;
wire R3C25_GT00;
wire R4C26_GB50;
wire R10C34_W10;
wire R18C4_GT00;
wire R22C39_GB30;
wire R10C28_W24;
wire R26C11_GBO0;
wire R15C1_GBO1;
wire R24C11_GB00;
wire R3C21_GB10;
wire R1C28_EW20;
wire R28C46_A6;
wire R12C24_GB50;
wire R14C40_GB20;
wire R14C45_GB30;
wire R26C32_GB60;
wire R6C8_GB20;
wire R26C23_GB00;
wire R28C7_C3;
wire R13C9_GB00;
wire R1C28_SEL7;
wire R4C21_GB20;
wire R9C30_GBO0;
wire R7C17_GB20;
wire R2C41_GB40;
wire R10C19_C2;
wire R28C25_N80;
wire R15C7_GB60;
wire R28C31_W26;
wire R11C38_GBO1;
wire R25C11_GB00;
wire R3C25_GBO1;
wire R7C11_GB40;
wire R28C28_B1;
wire R27C18_GBO0;
wire R28C7_W26;
wire R8C13_GB10;
wire R7C13_GB40;
wire R17C12_GB20;
wire R20C42_GB50;
wire R10C43_W11;
wire R28C13_SEL7;
wire R26C25_GT10;
wire R20C14_GB50;
wire R28C25_E80;
wire R12C8_GB60;
wire R28C22_CE1;
wire R23C12_GB50;
wire R16C44_GB20;
wire R5C22_GB50;
wire R15C13_GB60;
wire R17C29_GT00;
wire R9C33_GT00;
wire R2C23_GB10;
wire R7C40_GBO0;
wire R2C8_SPINE12;
wire R21C33_GB40;
wire R10C29_A5;
wire R28C7_Q1;
wire R16C21_GB30;
wire R1C47_E23;
wire R14C30_GB70;
wire R29C28_N13;
wire R12C3_GBO1;
wire R28C25_Q0;
wire R25C19_GB40;
wire R10C10_F4;
wire R9C12_GBO0;
wire R5C35_GB10;
wire R13C23_GB60;
wire R7C41_GB20;
wire R26C38_GBO1;
wire R15C41_GBO1;
wire R10C34_S80;
wire R28C19_SEL1;
wire R28C46_C2;
wire R20C36_GB50;
wire R28C40_B0;
wire R8C3_GT10;
wire R16C7_GBO0;
wire R8C46_GB60;
wire R13C20_GB50;
wire R20C46_GB20;
wire R4C27_GB10;
wire R25C17_GT10;
wire R6C39_GB20;
wire R14C45_GBO1;
wire R20C25_GB50;
wire R8C7_GB50;
wire R25C30_GB20;
wire R25C34_GB70;
wire R11C30_GB60;
wire R16C10_GT00;
wire R4C37_GBO0;
wire R5C31_GB60;
wire R10C37_S25;
wire R15C8_GB60;
wire R12C24_GBO0;
wire R17C25_GBO1;
wire R23C33_GT00;
wire R25C3_GBO0;
wire R10C10_Q1;
wire R2C26_SPINE10;
wire R9C46_GBO1;
wire R22C32_GB50;
wire R23C37_GB00;
wire R22C12_GB70;
wire R18C43_GB60;
wire R10C13_X01;
wire R28C22_Q5;
wire R13C37_GB60;
wire R28C13_S25;
wire R22C18_GB10;
wire R10C31_S80;
wire R25C28_GB60;
wire R17C15_GB30;
wire R24C8_GBO0;
wire R2C2_GBO0;
wire R28C4_W80;
wire R10C25_C2;
wire R24C35_GB10;
wire R28C34_B2;
wire R16C30_GBO1;
wire R10C37_D2;
wire R15C5_GB20;
wire R8C19_GB70;
wire R22C38_GBO1;
wire R24C20_GBO1;
wire R28C40_N22;
wire R9C5_GB50;
wire R25C35_GBO1;
wire R28C28_W23;
wire R10C19_W80;
wire R25C44_GB20;
wire R10C30_W27;
wire R10C26_E21;
wire R10C16_Q6;
wire R21C3_GB00;
wire R28C16_SN20;
wire R21C15_GB10;
wire R29C28_E83;
wire R22C29_GB10;
wire R3C3_GB00;
wire R9C20_GB10;
wire R21C5_GT00;
wire R16C4_GB10;
wire R4C26_GB20;
wire R17C15_GB60;
wire R24C9_GT00;
wire R26C12_GT10;
wire R21C21_GB50;
wire R18C11_GT00;
wire R28C7_S11;
wire R28C4_W82;
wire R6C10_GB60;
wire R11C19_GB70;
wire R22C18_GB30;
wire R6C45_GT00;
wire R3C5_GB50;
wire R28C40_E81;
wire R24C12_GB20;
wire R15C28_GB60;
wire R28C4_S11;
wire R28C7_Q6;
wire R10C30_UNK128;
wire R28C16_E21;
wire R24C45_GB70;
wire R6C40_GB30;
wire R6C44_GB10;
wire R10C43_S81;
wire R5C29_GB10;
wire R11C11_GBO1;
wire R13C22_GT10;
wire R11C2_GB30;
wire R18C30_GB40;
wire R7C11_GBO0;
wire R25C29_GB30;
wire R27C9_GT10;
wire R17C25_GT00;
wire R3C18_GBO1;
wire R13C8_GB50;
wire R10C28_C4;
wire R1C1_B2;
wire R9C34_GB10;
wire R20C33_GB70;
wire R28C22_B0;
wire R4C24_GB00;
wire R28C28_A3;
wire R28C31_S81;
wire R26C33_GT00;
wire R28C40_F0;
wire R9C6_GB20;
wire R6C10_GB40;
wire R10C13_E11;
wire R10C29_X07;
wire R5C29_GT00;
wire R2C38_GB50;
wire R16C33_GT10;
wire R10C26_SEL4;
wire R10C27_S13;
wire R2C8_GB70;
wire R10C26_X07;
wire R1C32_SEL7;
wire R26C24_GB10;
wire R22C44_GB30;
wire R12C39_GB60;
wire R17C42_GB70;
wire R11C40_GT10;
wire R9C28_GB60;
wire R13C30_GB70;
wire R10C16_LSR1;
wire R28C4_E82;
wire R11C21_GT00;
wire R21C3_GT10;
wire R8C1_GT00;
wire R28C25_SEL5;
wire R10C22_X03;
wire R28C16_F2;
wire R21C34_GT10;
wire R28C22_A5;
wire R14C17_GB00;
wire R26C4_GB70;
wire R7C44_GB20;
wire R17C35_GBO0;
wire R26C28_GB10;
wire R28C19_E24;
wire R28C40_A7;
wire R10C37_D3;
wire R28C37_N21;
wire R27C27_GB70;
wire R20C21_GB10;
wire R6C35_GT10;
wire R27C6_GBO1;
wire R25C44_GB30;
wire R18C14_GBO1;
wire R9C24_GB50;
wire R15C15_GB30;
wire R10C26_W23;
wire R2C19_GT10;
wire R28C13_A2;
wire R28C34_E13;
wire R26C17_GB50;
wire R16C35_GB10;
wire R28C28_N82;
wire R13C29_GT00;
wire R4C17_GB00;
wire R7C4_GB20;
wire R5C14_GB60;
wire R20C27_GB40;
wire R2C42_GB10;
wire R10C43_X03;
wire R29C28_C3;
wire R29C28_F7;
wire R10C30_E25;
wire R10C37_D1;
wire R11C36_GT10;
wire R1C28_X02;
wire R24C22_GB70;
wire R24C16_GBO1;
wire R27C40_GB20;
wire R25C20_GB50;
wire R10C22_SEL2;
wire R8C46_GT10;
wire R6C7_GB00;
wire R8C14_GB40;
wire R28C40_B7;
wire R14C14_GB50;
wire R7C6_GB00;
wire R26C38_GB70;
wire R10C7_A3;
wire R24C33_GB50;
wire R26C15_GB60;
wire R2C29_GB40;
wire R10C26_E24;
wire R10C37_Q0;
wire R18C22_GB30;
wire R18C16_GB30;
wire R18C24_GB50;
wire R22C41_GB60;
wire R28C22_W24;
wire R5C20_GB00;
wire R2C36_GB00;
wire R28C46_X05;
wire R10C40_E10;
wire R16C18_GBO1;
wire R4C43_GBO0;
wire R12C19_GT00;
wire R14C37_GB60;
wire R7C18_GB40;
wire R1C1_N83;
wire R28C7_SEL4;
wire R10C37_E82;
wire R16C10_GB30;
wire R17C34_GB40;
wire R16C11_GB70;
wire R12C1_GBO1;
wire R10C26_C5;
wire R6C37_GT10;
wire R27C27_GT10;
wire R3C25_GBO0;
wire R2C46_GB30;
wire R11C35_GB10;
wire R7C7_GBO1;
wire R3C16_GBO1;
wire R15C33_GBO1;
wire R10C16_W83;
wire R10C29_A6;
wire R28C10_S26;
wire R28C37_N23;
wire R25C6_GB70;
wire R7C34_GBO0;
wire R15C6_GB50;
wire R27C26_GB50;
wire R3C7_GB60;
wire R16C41_GB70;
wire R25C29_GB60;
wire R20C27_GT00;
wire R1C1_SEL1;
wire R24C1_GBO1;
wire R2C37_GB30;
wire R26C41_GBO1;
wire R28C40_CE0;
wire R10C28_B7;
wire R14C22_GB20;
wire R14C46_GB30;
wire R26C6_GT00;
wire R25C22_GB50;
wire R17C23_GB00;
wire R17C4_GB50;
wire R20C37_GB20;
wire R20C45_GB20;
wire R28C31_S26;
wire R17C44_GBO0;
wire R24C43_GT00;
wire R20C21_GB20;
wire R15C37_GB00;
wire R13C6_GBO1;
wire R18C40_GB10;
wire R21C42_GT00;
wire R10C19_D2;
wire R28C16_N83;
wire R25C23_GT00;
wire R28C46_B3;
wire R14C25_GB50;
wire R1C28_D0;
wire R28C37_Q0;
wire R5C10_GB60;
wire R20C27_GB50;
wire R17C46_GB70;
wire R10C31_E83;
wire R28C43_F5;
wire R28C25_Q2;
wire R10C10_S20;
wire R20C34_GB50;
wire R4C6_GT10;
wire R10C10_A5;
wire R10C10_A2;
wire R2C46_GB40;
wire R1C28_S83;
wire R8C21_GT10;
wire R10C7_W24;
wire R13C8_GBO0;
wire R10C25_SN20;
wire R29C28_CLK2;
wire R15C37_GB20;
wire R18C41_GB70;
wire R24C46_GB70;
wire R3C21_GB00;
wire R26C11_GB00;
wire R6C4_GB20;
wire R6C19_GB70;
wire R17C36_GB60;
wire R28C31_F2;
wire R8C30_GB60;
wire R9C26_GB10;
wire R17C46_GT10;
wire R24C26_GB10;
wire R9C18_GB10;
wire R25C2_GBO0;
wire R26C9_GB70;
wire R10C30_W25;
wire R16C4_GB00;
wire R5C42_GB60;
wire R28C22_C2;
wire R10C34_X07;
wire R3C17_GB30;
wire R16C39_GT00;
wire R2C3_GB60;
wire R20C26_GB10;
wire R20C46_SPINE26;
wire R13C7_GBO1;
wire R10C10_F5;
wire R28C13_E80;
wire R28C16_F7;
wire R28C22_D7;
wire R2C2_GB60;
wire R25C23_GB40;
wire R6C7_GT10;
wire R13C21_GB00;
wire R4C40_GB70;
wire R17C38_GBO0;
wire R10C19_A0;
wire R13C7_GB40;
wire R16C11_GB50;
wire R15C6_GB10;
wire R28C34_LSR1;
wire R27C22_GBO0;
wire R10C40_E80;
wire R28C28_Q1;
wire R3C35_GB50;
wire R28C31_E27;
wire R26C10_GB00;
wire R13C35_GB30;
wire R16C4_GB40;
wire R1C28_X04;
wire R23C44_GB70;
wire R10C40_EW10;
wire R17C39_GB20;
wire R4C29_GT10;
wire R16C31_GT00;
wire R10C7_F0;
wire R28C34_E80;
wire R8C21_GB30;
wire R10C25_B0;
wire R10C13_S20;
wire R9C16_GB60;
wire R26C2_GBO0;
wire R1C1_N24;
wire R26C41_GB20;
wire R5C42_GB10;
wire R10C29_C4;
wire R15C19_GBO0;
wire R27C39_GBO1;
wire R10C16_W12;
wire R22C36_GBO0;
wire R15C40_GB00;
wire R10C10_N13;
wire R17C20_GT00;
wire R4C32_GB40;
wire R28C25_LSR1;
wire R10C31_W27;
wire R6C13_GB10;
wire R28C19_A5;
wire R8C19_GBO1;
wire R16C9_GB50;
wire R22C17_GB00;
wire R27C16_GB30;
wire R13C15_GB40;
wire R16C27_GB30;
wire R26C15_GB20;
wire R10C25_C7;
wire R3C9_GB10;
wire R8C8_GBO1;
wire R28C40_A3;
wire R1C32_CLK0;
wire R24C27_GB50;
wire R8C33_GB20;
wire R3C25_GB40;
wire R28C19_N12;
wire R16C25_GB60;
wire R27C18_GB70;
wire R28C22_W26;
wire R13C18_GB70;
wire R21C29_GB20;
wire R10C25_F1;
wire R17C34_GT00;
wire R20C27_SPINE21;
wire R16C21_GBO0;
wire R23C8_GBO1;
wire R22C46_GB30;
wire R10C30_S10;
wire R20C1_GT10;
wire R16C12_GT10;
wire R4C21_GB00;
wire R5C21_GB60;
wire R18C35_GB00;
wire R22C30_GBO0;
wire R4C18_GB70;
wire R27C14_GB30;
wire R20C33_GBO1;
wire R9C38_GB20;
wire R28C25_SEL4;
wire R18C27_GB00;
wire R24C14_GB20;
wire R10C34_N13;
wire R7C34_GB00;
wire R21C10_GB60;
wire R10C28_EW10;
wire R28C43_X01;
wire R7C20_GBO1;
wire R28C7_S83;
wire R24C8_GB60;
wire R16C26_GT10;
wire R13C34_GT00;
wire R24C26_GB30;
wire R7C15_GBO1;
wire R12C3_GB10;
wire R10C19_W82;
wire R4C2_GB10;
wire R5C27_GBO0;
wire R20C4_GB30;
wire R28C7_CE2;
wire R28C16_N20;
wire R2C5_GB60;
wire R16C36_GB10;
wire R10C27_E13;
wire R24C3_GBO1;
wire R10C10_X05;
wire R29C28_W24;
wire R14C35_GT00;
wire R28C19_N27;
wire R27C17_GB50;
wire R17C36_GT00;
wire R18C37_GB00;
wire R28C16_A2;
wire R10C40_W25;
wire R25C21_GB40;
wire R11C11_GBO0;
wire R16C20_GB60;
wire R24C20_GB20;
wire R12C30_GB10;
wire R6C39_GB40;
wire R5C46_GB10;
wire R4C27_GB30;
wire R24C46_GT10;
wire R7C2_GB30;
wire R22C3_GT10;
wire R3C15_GB60;
wire R24C4_GB10;
wire R21C12_GB40;
wire R11C20_GB40;
wire R7C36_GBO1;
wire R16C33_GB40;
wire R25C40_GBO1;
wire R15C4_GB50;
wire R10C10_Q4;
wire R10C26_S12;
wire R27C31_GB00;
wire R25C16_GT10;
wire R24C12_GB40;
wire R22C31_GB30;
wire R22C19_GB10;
wire R27C30_GT00;
wire R15C31_GB20;
wire R15C43_GBO0;
wire R10C37_D4;
wire R15C14_GB30;
wire R28C4_A3;
wire R28C34_E12;
wire R28C34_N81;
wire R24C38_GB10;
wire R27C10_GB50;
wire R5C14_GB20;
wire R26C34_GT00;
wire R7C34_GB70;
wire R12C24_GB60;
wire R28C31_W20;
wire R28C19_N25;
wire R20C10_GB30;
wire R21C22_GB20;
wire R3C28_GB10;
wire R20C45_GB00;
wire R13C24_GB50;
wire R28C19_S82;
wire R7C10_GB10;
wire R11C9_GB10;
wire R2C40_GB40;
wire R15C29_GB60;
wire R10C29_SEL3;
wire R7C12_GB30;
wire R25C16_GBO0;
wire R23C35_GB70;
wire R10C29_C3;
wire R8C23_GBO0;
wire R2C26_GB30;
wire R24C10_GB20;
wire R17C28_GT00;
wire R25C40_GT00;
wire R14C25_GBO0;
wire R15C26_GB70;
wire R5C20_GB60;
wire R11C24_GB00;
wire R12C26_GBO0;
wire R24C25_GT10;
wire R13C46_GT10;
wire R23C23_GB20;
wire R22C34_GT10;
wire R25C13_GT00;
wire R20C26_GB20;
wire R23C4_GB30;
wire R23C15_GB70;
wire R5C12_GB40;
wire R4C11_GB00;
wire R4C26_GB30;
wire R24C21_GB00;
wire R10C22_W81;
wire R10C37_W26;
wire R1C28_E23;
wire R26C43_GB50;
wire R28C25_N10;
wire R27C46_GBO0;
wire R10C16_E27;
wire R23C30_GB40;
wire R24C19_GB20;
wire R12C7_GT00;
wire R28C16_N11;
wire R23C38_GB70;
wire R25C19_GB10;
wire R10C22_S13;
wire R4C38_GB30;
wire R13C31_GB60;
wire R10C25_W82;
wire R2C4_SPINE12;
wire R28C10_N27;
wire R23C34_GB30;
wire R28C7_F4;
wire R10C37_N20;
wire R25C24_GB70;
wire R29C28_B3;
wire R23C8_GT00;
wire R9C25_GB50;
wire R4C12_GBO1;
wire R3C43_GT10;
wire R1C1_D0;
wire R26C37_GB30;
wire R16C15_GB70;
wire R16C2_GB50;
wire R22C6_GB10;
wire R8C14_GBO0;
wire R24C5_GB20;
wire R3C19_GB70;
wire R10C19_D4;
wire R5C33_GB40;
wire R2C43_GB10;
wire R13C30_GB20;
wire R6C12_GB40;
wire R1C47_W80;
wire R5C30_GB40;
wire R1C28_S11;
wire R25C14_GT10;
wire R10C37_CLK1;
wire R13C11_GB40;
wire R3C24_GB30;
wire R7C27_GB40;
wire R22C21_GB00;
wire R21C15_GBO1;
wire R7C18_GB10;
wire R28C31_Q6;
wire R1C47_X03;
wire R10C30_W24;
wire R28C37_Q6;
wire R7C11_GB70;
wire R7C14_GB40;
wire R28C28_F5;
wire R3C18_GB30;
wire R8C21_GB00;
wire R2C8_GT00;
wire R14C13_GBO0;
wire R17C29_GBO1;
wire R12C33_GB10;
wire R25C2_GB10;
wire R28C46_W27;
wire R6C36_GB50;
wire R13C18_GT00;
wire R10C29_S21;
wire R10C10_D1;
wire R22C35_GB00;
wire R12C39_GB40;
wire R10C25_LSR2;
wire R12C35_GT10;
wire R10C27_F3;
wire R17C6_GB70;
wire R11C13_GT10;
wire R7C36_GB50;
wire R4C36_GT00;
wire R10C16_A1;
wire R15C42_GT10;
wire R21C5_GT10;
wire R3C26_GB10;
wire R27C38_GT00;
wire R10C7_F6;
wire R15C39_GB30;
wire R14C18_GT00;
wire R10C25_N22;
wire R3C6_GB20;
wire R28C22_N27;
wire R15C11_GBO1;
wire R28C22_N11;
wire R18C26_GB20;
wire R28C40_W13;
wire R5C10_GBO0;
wire R13C45_GB10;
wire R28C16_SEL5;
wire R28C28_N10;
wire R22C34_GBO1;
wire R3C5_GB40;
wire R21C13_GB70;
wire R13C33_GB30;
wire R23C24_GB00;
wire R28C40_SEL6;
wire R14C24_GB20;
wire R2C13_SPINE11;
wire R7C21_GB20;
wire R23C8_GB20;
wire R14C1_GBO1;
wire R6C41_GB50;
wire R15C23_GB10;
wire R1C28_B5;
wire R13C33_GT10;
wire R10C31_C5;
wire R13C35_GB50;
wire R18C42_GB60;
wire R9C22_GB50;
wire R18C16_GB70;
wire R22C5_GB30;
wire R22C15_GB20;
wire R10C19_N27;
wire R26C21_GB10;
wire R20C32_GBO0;
wire R7C26_GBO0;
wire R17C42_GB30;
wire R17C31_GBO0;
wire R10C19_N21;
wire R10C22_E20;
wire R10C34_B7;
wire R11C8_GBO0;
wire R9C23_GBO1;
wire R20C7_GB60;
wire R12C36_GB40;
wire R11C44_GB40;
wire R28C19_F3;
wire R10C43_A5;
wire R17C9_GB30;
wire R25C36_GB00;
wire R11C12_GB10;
wire R22C45_GB20;
wire R13C34_GB30;
wire R7C15_GB10;
wire R7C13_GB00;
wire R4C16_GB00;
wire R17C13_GB60;
wire R10C31_W23;
wire R27C7_GBO0;
wire R27C9_GT00;
wire R25C33_GBO1;
wire R4C3_GB30;
wire R1C32_E10;
wire R28C34_S22;
wire R14C35_GB20;
wire R10C29_UNK128;
wire R21C18_GB40;
wire R15C22_GB00;
wire R10C37_N21;
wire R27C41_GBO1;
wire R23C39_GBO0;
wire R10C13_EW10;
wire R16C15_GB20;
wire R22C26_GBO1;
wire R28C19_W24;
wire R27C30_GB10;
wire R6C24_GT00;
wire R11C44_GB20;
wire R10C43_EW10;
wire R28C10_F4;
wire R28C28_B3;
wire R22C38_GT10;
wire R17C21_GB40;
wire R25C39_GBO1;
wire R4C9_GB20;
wire R12C44_GB60;
wire R10C37_B3;
wire R2C17_GT00;
wire R16C2_GB00;
wire R12C43_GB10;
wire R20C41_GB70;
wire R24C24_GB30;
wire R23C46_GBO0;
wire R27C46_GB20;
wire R10C7_W26;
wire R4C36_GT10;
wire R7C36_GT10;
wire R4C14_GB10;
wire R5C3_GB10;
wire R11C12_GBO0;
wire R9C11_GB30;
wire R8C20_GB70;
wire R26C42_GB10;
wire R12C4_GT00;
wire R25C6_GB10;
wire R10C37_X03;
wire R28C7_E81;
wire R4C24_GB60;
wire R28C10_F1;
wire R25C24_GB60;
wire R22C4_GB20;
wire R12C25_GBO1;
wire R11C38_GB50;
wire R21C33_GBO1;
wire R1C47_E13;
wire R10C7_W11;
wire R26C3_GT00;
wire R23C14_GB00;
wire R10C40_N27;
wire R7C3_GB20;
wire R28C7_SN20;
wire R20C20_GT00;
wire R15C34_GT10;
wire R4C10_GB10;
wire R21C15_GB40;
wire R27C27_GBO1;
wire R15C16_GB60;
wire R13C26_GB70;
wire R28C46_N27;
wire R15C24_GB60;
wire R8C18_GB10;
wire R17C40_GBO1;
wire R28C43_W23;
wire R15C7_GB30;
wire R28C13_E21;
wire R20C32_GB50;
wire R27C34_GB30;
wire R29C28_F4;
wire R25C35_GB10;
wire R13C41_GB70;
wire R29C28_Q3;
wire R1C47_D6;
wire R28C16_D1;
wire R15C8_GB30;
wire R16C34_GBO0;
wire R9C32_GB10;
wire R20C18_GB10;
wire R25C23_GT10;
wire R12C21_GB70;
wire R9C27_GB70;
wire R3C30_GB70;
wire R9C4_GB10;
wire R21C44_GT00;
wire R23C37_GBO1;
wire R28C28_N20;
wire R24C41_GB70;
wire R8C23_GB40;
wire R14C5_GB30;
wire R3C36_GB70;
wire R14C43_GB20;
wire R25C7_GB10;
wire R10C40_S10;
wire R28C25_W81;
wire R10C40_F5;
wire R10C28_F5;
wire R18C31_GB40;
wire R10C26_E11;
wire R10C43_Q3;
wire R24C37_GBO0;
wire R11C42_GT10;
wire R21C1_GT10;
wire R18C32_GT10;
wire R25C41_GBO0;
wire R10C29_W21;
wire R28C25_C6;
wire R16C20_GB50;
wire R9C39_GBO0;
wire R28C34_S26;
wire R28C10_S11;
wire R26C4_GB50;
wire R12C29_GBO0;
wire R28C13_LSR0;
wire R3C25_GB50;
wire R18C5_GB20;
wire R10C37_EW20;
wire R1C32_N23;
wire R28C22_SEL1;
wire R2C35_GB60;
wire R14C7_GB50;
wire R12C9_GB60;
wire R17C31_GB00;
wire R16C37_GB70;
wire R1C32_N13;
wire R10C43_F1;
wire R4C46_GT10;
wire R21C40_GB10;
wire R13C33_GBO0;
wire R10C25_S11;
wire R7C19_GBO1;
wire R12C33_GB40;
wire R20C11_GB00;
wire R21C8_GT10;
wire R28C16_F3;
wire R20C13_GT00;
wire R10C30_CE2;
wire R28C16_X02;
wire R18C3_GBO0;
wire R11C36_GB40;
wire R21C17_GB60;
wire R15C27_GB00;
wire R23C8_GB00;
wire R11C19_GB00;
wire R18C2_GB50;
wire R18C21_GB60;
wire R20C16_GB30;
wire R6C30_GBO0;
wire R21C46_GB20;
wire R18C32_GB60;
wire R11C20_GB00;
wire R8C36_GB00;
wire R10C43_N81;
wire R12C5_GB00;
wire R27C14_GB10;
wire R3C41_GB60;
wire R7C23_GB20;
wire R1C32_A5;
wire R26C18_GB40;
wire R16C27_GT10;
wire R8C25_GT00;
wire R4C8_GB60;
wire R25C10_GB10;
wire R20C4_GBO0;
wire R2C26_GBO0;
wire R12C18_GB20;
wire R22C42_GB30;
wire R26C35_GB70;
wire R2C24_GBO0;
wire R10C25_N80;
wire R10C19_N20;
wire R15C27_GT10;
wire R16C34_GB20;
wire R13C36_GB50;
wire R16C8_GT00;
wire R2C14_GBO1;
wire R12C40_GT10;
wire R26C13_GT10;
wire R21C12_GB60;
wire R26C16_GB40;
wire R14C16_GB60;
wire R28C4_S21;
wire R14C6_GB20;
wire R28C10_SEL3;
wire R1C47_N12;
wire R10C37_S81;
wire R16C23_GBO0;
wire R12C25_GB10;
wire R28C37_X03;
wire R12C46_GB10;
wire R8C17_GB70;
wire R10C25_B1;
wire R24C17_GB00;
wire R23C28_GB30;
wire R24C27_GBO1;
wire R2C11_SPINE13;
wire R25C17_GB50;
wire R22C9_GT00;
wire R27C21_GB60;
wire R6C8_GBO0;
wire R25C14_GB60;
wire R4C42_GB20;
wire R25C3_GB30;
wire R1C47_A2;
wire R16C16_GBO1;
wire R1C32_S26;
wire R10C16_S24;
wire R20C8_GB00;
wire R9C1_GBO1;
wire R8C33_GT00;
wire R24C26_GB00;
wire R28C28_X03;
wire R8C23_GB70;
wire R29C28_X07;
wire R17C37_GB00;
wire R7C38_GB00;
wire R28C19_W22;
wire R7C10_GB30;
wire R23C2_GB70;
wire R26C39_GT10;
wire R25C3_GB70;
wire R20C15_GB20;
wire R4C2_GT10;
wire R7C46_GB10;
wire R1C32_E21;
wire R10C27_B0;
wire R25C46_GT10;
wire R10C13_C3;
wire R10C16_S13;
wire R16C31_GT10;
wire R26C10_GB50;
wire R28C25_F3;
wire R27C31_GT10;
wire R27C39_GB60;
wire R4C10_GT10;
wire R11C13_GB50;
wire R14C13_GBO1;
wire R6C10_GT10;
wire R21C14_GB10;
wire R11C33_GB30;
wire R5C45_GB60;
wire R10C10_N27;
wire R10C13_CLK2;
wire R10C26_CLK0;
wire R28C25_S20;
wire R17C14_GT00;
wire R4C29_GBO1;
wire R28C40_C0;
wire R5C13_GB50;
wire R1C32_Q0;
wire R3C42_GT10;
wire R28C7_Q7;
wire R17C44_GT00;
wire R28C46_N25;
wire R4C32_GB10;
wire R28C46_F3;
wire R8C18_GB20;
wire R28C31_X06;
wire R14C42_GB50;
wire R28C46_SEL4;
wire R2C16_GB70;
wire R2C44_GB60;
wire R24C33_GB00;
wire R28C4_X05;
wire R28C7_W11;
wire R21C39_GB40;
wire R24C39_GBO1;
wire R10C27_A0;
wire R1C1_Q2;
wire R26C42_GB40;
wire R8C15_GB70;
wire R4C33_GB10;
wire R1C28_N11;
wire R28C46_F4;
wire R2C9_GB20;
wire R4C24_GB30;
wire R4C9_GT00;
wire R22C27_GB60;
wire R10C30_E10;
wire R28C40_CE1;
wire R10C7_W12;
wire R6C41_GB40;
wire R26C13_GT00;
wire R5C23_GB10;
wire R10C22_CE0;
wire R10C22_Q7;
wire R5C35_GB00;
wire R12C27_GBO1;
wire R24C42_GBO0;
wire R25C41_GB70;
wire R13C2_GBO0;
wire R23C41_GT00;
wire R11C40_GT00;
wire R27C22_GB00;
wire R28C22_N81;
wire R17C3_GB70;
wire R10C31_N27;
wire R28C22_A2;
wire R18C19_GB10;
wire R10C40_D7;
wire R28C10_N23;
wire R14C20_GB00;
wire R15C38_GBO1;
wire R3C45_GB50;
wire R7C42_GB50;
wire R29C28_B6;
wire R10C28_UNK126;
wire R28C43_W21;
wire R3C40_GB40;
wire R8C26_GT10;
wire R14C13_GT10;
wire R6C17_GBO0;
wire R10C19_A3;
wire R28C28_S22;
wire R10C10_C3;
wire R10C37_F5;
wire R13C23_GB00;
wire R15C31_GB30;
wire R21C43_GB40;
wire R10C27_SEL0;
wire R25C24_GB10;
wire R10C16_N12;
wire R10C7_SN20;
wire R28C19_A7;
wire R26C46_GT00;
wire R25C44_GBO1;
wire R21C23_GB00;
wire R8C12_GB10;
wire R2C24_GB50;
wire R5C26_GT00;
wire R16C28_GB20;
wire R25C42_GBO1;
wire R26C43_GB00;
wire R5C27_GB20;
wire R28C28_N24;
wire R13C33_GT00;
wire R22C31_GB40;
wire R7C6_GBO0;
wire R10C26_SEL5;
wire R12C32_GB20;
wire R3C6_GB30;
wire R25C4_GB00;
wire R15C26_GB60;
wire R9C31_GB00;
wire R6C38_GB20;
wire R2C38_GB30;
wire R8C39_GBO1;
wire R16C40_GBO1;
wire R23C3_GB40;
wire R10C26_F6;
wire R10C28_B6;
wire R10C43_SEL0;
wire R13C18_GB00;
wire R10C16_SN10;
wire R4C41_GB30;
wire R5C31_GB10;
wire R4C31_GT00;
wire R17C33_GB00;
wire R10C31_D0;
wire R10C40_E25;
wire R28C31_W22;
wire R12C8_GBO0;
wire R27C7_GT10;
wire R24C44_GT10;
wire R28C7_X08;
wire R24C24_GT00;
wire R10C29_B2;
wire R25C12_GB00;
wire R26C26_GB40;
wire R9C19_GB10;
wire R28C28_SEL5;
wire R8C10_GB70;
wire R13C4_GB70;
wire R4C28_GT10;
wire R3C11_GBO1;
wire R24C37_GB00;
wire R8C18_GT00;
wire R12C33_GB70;
wire R10C25_Q3;
wire R5C20_GB50;
wire R16C4_GB20;
wire R10C30_W26;
wire R14C38_GBO0;
wire R10C26_B6;
wire R4C40_GB30;
wire R8C4_GB50;
wire R28C25_S81;
wire R24C29_GBO0;
wire R25C32_GB50;
wire R18C18_GB50;
wire R10C30_Q6;
wire R3C38_GB00;
wire R12C11_GB40;
wire R10C31_X04;
wire R2C27_GT10;
wire R10C26_S22;
wire R13C28_GT00;
wire R10C29_Q2;
wire R20C34_GT00;
wire R28C10_C7;
wire R23C46_GB30;
wire R22C14_GT00;
wire R11C7_GT10;
wire R10C34_W12;
wire R23C40_GB30;
wire R2C42_GB30;
wire R28C28_W13;
wire R10C22_B1;
wire R23C34_GT00;
wire R26C38_GT10;
wire R1C28_N21;
wire R18C23_GBO1;
wire R4C43_GB70;
wire R7C28_GB20;
wire R2C16_SPINE8;
wire R4C31_GT10;
wire R14C16_GB30;
wire R26C9_GB40;
wire R6C46_GBO0;
wire R10C10_C5;
wire R10C31_B6;
wire R10C34_F3;
wire R28C22_B2;
wire R17C38_GB20;
wire R28C28_A7;
wire R22C13_GB70;
wire R21C30_GB00;
wire R24C5_GB50;
wire R22C46_GB10;
wire R17C17_GB40;
wire R21C10_GBO1;
wire R16C41_GBO0;
wire R21C28_GB40;
wire R12C28_GB60;
wire R2C37_GB10;
wire R22C44_GB10;
wire R15C25_GB50;
wire R28C46_SEL3;
wire R20C44_GB50;
wire R28C37_E26;
wire R8C6_GB30;
wire R14C40_GBO0;
wire R20C45_SPINE27;
wire R10C25_CLK2;
wire R3C40_GB60;
wire R9C16_GT00;
wire R10C43_F7;
wire R11C10_GT10;
wire R27C46_GT10;
wire R27C40_GB00;
wire R2C38_GB20;
wire R24C44_GB70;
wire R4C46_GB10;
wire R6C23_GB70;
wire R17C30_GB40;
wire VCC;
wire R20C29_GB30;
wire R16C29_GB10;
wire R20C17_GB70;
wire R12C27_GB50;
wire R7C33_GB60;
wire R10C34_Q5;
wire R28C25_Q1;
wire R23C27_GT10;
wire R1C28_W23;
wire R1C28_E11;
wire R10C28_CLK1;
wire R28C13_X01;
wire R14C4_GB60;
wire R9C6_GB30;
wire R27C15_GB60;
wire R16C26_GB50;
wire R4C25_GBO0;
wire R26C39_GB50;
wire R25C33_GT10;
wire R9C27_GB00;
wire R2C31_SPINE1;
wire R17C33_GT00;
wire R6C6_GB20;
wire R3C19_GB60;
wire R5C34_GB30;
wire R10C30_N20;
wire R28C40_N23;
wire R10C34_N11;
wire R28C31_B5;
wire R18C28_GB30;
wire R11C40_GB20;
wire R18C5_GB30;
wire R10C10_W83;
wire R4C22_GB30;
wire R17C3_GB50;
wire R7C22_GBO1;
wire R21C29_GB10;
wire R20C17_GB30;
wire R23C17_GB30;
wire R28C46_W20;
wire R4C27_GT00;
wire R10C22_X06;
wire R22C39_GB20;
wire R15C12_GB00;
wire R17C19_GB00;
wire R15C9_GBO0;
wire R26C12_GBO1;
wire R27C19_GT00;
wire R15C28_GB10;
wire R17C26_GB00;
wire R17C11_GB50;
wire R5C43_GB00;
wire R22C2_GB50;
wire R1C28_CE0;
wire R17C11_GBO1;
wire R5C8_GB00;
wire R11C38_GBO0;
wire R25C45_GB60;
wire R12C6_GT10;
wire R7C45_GB40;
wire R28C40_SEL0;
wire R13C18_GT10;
wire R12C20_GB60;
wire R6C44_GB30;
wire R10C25_CLK1;
wire R10C43_CE1;
wire R18C21_GBO0;
wire R1C32_S21;
wire R3C12_GB20;
wire R21C26_GB60;
wire R2C43_GB00;
wire R2C25_GB40;
wire R11C6_GB70;
wire R2C25_GBO1;
wire R18C2_GT10;
wire R28C31_X08;
wire R10C19_E80;
wire R15C17_GBO0;
wire R12C44_GB20;
wire R28C13_N22;
wire R18C44_GB70;
wire R17C44_GB30;
wire R9C46_GB40;
wire R8C45_GT10;
wire R8C10_GT00;
wire R6C12_GB20;
wire R28C4_A4;
wire R28C7_X06;
wire R10C22_SN10;
wire R12C14_GB30;
wire R28C37_S25;
wire R21C36_GB50;
wire R12C28_GB40;
wire R13C37_GB50;
wire R18C32_GB40;
wire R9C42_GB70;
wire R15C44_GB50;
wire R10C13_X04;
wire R28C13_A4;
wire R25C3_GT00;
wire R7C34_GT00;
wire R28C19_SEL0;
wire R26C23_GBO1;
wire R26C10_GB30;
wire R21C40_GB30;
wire R3C43_GB70;
wire R28C25_S24;
wire R3C13_GB10;
wire R2C40_SPINE4;
wire R11C10_GB40;
wire R4C18_GT00;
wire R6C11_GBO1;
wire R2C18_GB60;
wire R21C12_GB00;
wire R18C46_GBO1;
wire R11C19_GB20;
wire R4C4_GBO0;
wire R20C25_GT10;
wire R21C15_GB00;
wire R24C35_GB00;
wire R20C39_GBO0;
wire R10C16_C5;
wire R18C33_GT00;
wire R11C42_GB40;
wire R2C19_GBO1;
wire R20C21_GB40;
wire R28C16_N26;
wire R9C7_GB30;
wire R16C9_GB30;
wire R16C2_GB40;
wire R24C7_GB20;
wire R8C45_GB50;
wire R10C10_EW10;
wire R13C4_GBO0;
wire R12C6_GB60;
wire R8C42_GBO1;
wire R28C7_N13;
wire R28C37_F5;
wire R27C19_GB30;
wire R9C15_GB30;
wire R24C18_GB20;
wire R27C4_GB70;
wire R28C28_C4;
wire R4C16_GBO1;
wire R7C14_GB10;
wire R6C28_GB40;
wire R14C5_GB20;
wire R10C30_X05;
wire R24C18_GBO0;
wire R28C13_S22;
wire R26C11_GT00;
wire R10C28_W26;
wire R10C7_F7;
wire R28C43_X04;
wire R14C7_GT10;
wire R20C41_GB60;
wire R4C19_GB10;
wire R22C35_GB60;
wire R7C29_GB20;
wire R11C18_GB50;
wire R15C46_GB60;
wire R28C16_N22;
wire R28C13_F7;
wire R24C39_GB40;
wire R10C29_D0;
wire R27C38_GB00;
wire R14C10_GB70;
wire R17C39_GBO1;
wire R28C34_W25;
wire R24C14_GBO1;
wire R27C12_GT00;
wire R25C22_GB70;
wire R27C43_GB50;
wire R26C27_GBO1;
wire R24C23_GT00;
wire R23C30_GT10;
wire R11C15_GB40;
wire R24C41_GB20;
wire R13C26_GB20;
wire R26C31_GB50;
wire R4C41_GB60;
wire R17C24_GBO1;
wire R4C12_GB60;
wire R18C13_GB70;
wire R23C42_GB00;
wire R20C40_GB20;
wire R22C38_GB30;
wire R18C30_GB70;
wire R1C47_C3;
wire R25C37_GB60;
wire R10C16_SEL3;
wire R6C38_GB50;
wire R11C31_GB30;
wire R26C33_GBO1;
wire R10C25_W21;
wire R8C26_GBO0;
wire R6C24_GB50;
wire R10C22_A7;
wire R13C9_GBO1;
wire R9C21_GB70;
wire R9C45_GB00;
wire R5C22_GBO1;
wire R16C40_GT10;
wire R22C8_GB30;
wire R18C29_GB30;
wire R5C10_GB30;
wire R28C7_N27;
wire R10C10_A3;
wire R6C26_GT00;
wire R4C17_GB50;
wire R23C24_GB50;
wire R20C10_GBO1;
wire R2C45_GB60;
wire R11C30_GB00;
wire R10C30_SPINE4;
wire R17C26_GB30;
wire R8C8_GB30;
wire R25C36_GB10;
wire R22C35_GB20;
wire R23C6_GB00;
wire R12C26_GBO1;
wire R18C37_GB10;
wire R10C22_Q5;
wire R28C13_D3;
wire R10C16_W22;
wire R12C21_GB10;
wire R9C18_GB50;
wire R17C31_GB20;
wire R14C4_GBO0;
wire R13C6_GB60;
wire R1C47_W26;
wire R10C16_E13;
wire R5C24_GT10;
wire R24C9_GB30;
wire R28C40_D0;
wire R20C36_GB10;
wire R3C38_GB70;
wire R5C10_GB20;
wire R24C18_GB00;
wire R18C7_GBO0;
wire R13C12_GB10;
wire R27C14_GT10;
wire R10C28_X08;
wire R14C19_GB50;
wire R28C22_W20;
wire R4C28_GT00;
wire R7C16_GB00;
wire R9C36_GBO1;
wire R8C46_GB40;
wire R28C4_W81;
wire R6C27_GB10;
wire R28C16_LSR2;
wire R15C31_GBO1;
wire R9C6_GT10;
wire R11C25_GB60;
wire R22C7_GB30;
wire R15C27_GB70;
wire R12C13_GB30;
wire R2C3_SPINE9;
wire R25C31_GT10;
wire R4C35_GBO1;
wire R26C45_GBO0;
wire R10C43_S80;
wire R28C28_S24;
wire R28C43_N21;
wire R7C45_GT10;
wire R7C20_GBO0;
wire R28C22_X05;
wire R27C22_GB40;
wire R29C28_CLK0;
wire R26C29_GB10;
wire R16C37_GB40;
wire R28C7_A7;
wire R13C46_GB20;
wire R27C40_GT10;
wire R10C13_N82;
wire R28C46_X03;
wire R10C19_S83;
wire R27C5_GB50;
wire R10C26_X02;
wire R17C17_GB20;
wire R4C33_GB60;
wire R16C14_GT10;
wire R11C30_GT00;
wire R6C43_GT10;
wire R24C34_GB30;
wire R10C28_E12;
wire R24C28_GB10;
wire R11C17_GBO1;
wire R25C22_GBO0;
wire R24C37_GB20;
wire R7C14_GB00;
wire R1C28_N12;
wire R17C13_GB20;
wire R17C20_GB40;
wire R24C22_GB00;
wire R10C13_B0;
wire R16C27_GB40;
wire R22C21_GB10;
wire R20C26_GB50;
wire R25C28_GB10;
wire R4C31_GB50;
wire R15C33_GBO0;
wire R10C34_N23;
wire R12C23_GT00;
wire R2C41_GT10;
wire R28C46_E21;
wire R28C34_A3;
wire R28C40_E82;
wire R10C40_SEL2;
wire R6C17_GBO1;
wire R9C6_GB60;
wire R28C25_B3;
wire R2C38_GT00;
wire R11C10_GB00;
wire R23C39_GB00;
wire R21C36_GBO1;
wire R26C11_GT10;
wire R20C40_GB70;
wire R18C31_GB30;
wire R10C26_CE0;
wire R24C44_GB00;
wire R8C3_GB60;
wire R4C18_GB60;
wire R20C43_GT10;
wire R23C35_GB40;
wire R29C28_F5;
wire R7C43_GB10;
wire R13C21_GB20;
wire R5C30_GB60;
wire R22C8_GB20;
wire R28C40_N21;
wire R28C40_SN20;
wire R22C43_GBO1;
wire R16C16_GB40;
wire R2C9_GBO0;
wire R11C14_GB40;
wire R10C43_CLK0;
wire R23C13_GT00;
wire R23C31_GB60;
wire R28C7_N25;
wire R7C39_GB00;
wire R10C13_SN20;
wire R28C4_EW10;
wire R11C5_GB60;
wire R21C17_GB30;
wire R28C43_E13;
wire R16C24_GBO1;
wire R8C37_GT00;
wire R12C37_GB40;
wire R9C12_GB00;
wire R28C34_A7;
wire R9C34_GB70;
wire R10C16_S22;
wire R15C6_GB40;
wire R18C19_GBO0;
wire R21C17_GT10;
wire R20C33_GT10;
wire R25C21_GB20;
wire R15C33_GB00;
wire R11C29_GB70;
wire R10C28_Q2;
wire R10C13_W80;
wire R10C34_C6;
wire R20C12_GB30;
wire R28C37_X06;
wire R20C32_GB20;
wire R20C11_GB40;
wire R11C31_GB60;
wire R4C24_GT00;
wire R26C37_GB20;
wire R23C41_GB50;
wire R10C13_Q1;
wire R10C31_B3;
wire R10C27_Q7;
wire R21C24_GB10;
wire R5C18_GB60;
wire R23C1_GBO0;
wire R10C31_SEL6;
wire R10C10_E82;
wire R11C28_GB50;
wire R10C10_N24;
wire R10C31_S24;
wire R28C37_Q3;
wire R1C28_E83;
wire R20C36_SPINE24;
wire R12C45_GT00;
wire R4C3_GB10;
wire R26C14_GB20;
wire R4C41_GT10;
wire R9C36_GB40;
wire R27C28_GB40;
wire R24C41_GB50;
wire R8C14_GB50;
wire R17C29_GB10;
wire R10C22_A1;
wire R5C5_GT00;
wire R10C28_W22;
wire R7C13_GT10;
wire R11C20_GBO0;
wire R20C46_GB40;
wire R3C11_GBO0;
wire R17C9_GT00;
wire R21C46_GBO1;
wire R28C25_D0;
wire R2C5_GB00;
wire R16C2_GT10;
wire R21C9_GB10;
wire R12C35_GB60;
wire R25C46_GB70;
wire R7C32_GB00;
wire R28C19_E83;
wire R13C32_GB30;
wire R11C24_GB30;
wire R5C1_GT10;
wire R28C4_X02;
wire R6C2_GBO1;
wire R2C24_GB60;
wire R1C1_W24;
wire R23C43_GB20;
wire R10C13_N25;
wire R10C22_Q2;
wire R10C25_S26;
wire R16C23_GT10;
wire R10C28_SN20;
wire R15C32_GT10;
wire R17C29_GB00;
wire R20C41_GBO1;
wire R25C30_GB30;
wire R12C42_GB50;
wire R20C37_GB30;
wire R28C37_X02;
wire R27C37_GBO1;
wire R25C5_GB00;
wire R9C27_GT00;
wire R20C22_GB70;
wire R26C41_GB40;
wire R1C32_SEL4;
wire R10C29_B4;
wire R15C39_GT00;
wire R5C16_GT10;
wire R2C40_GB30;
wire R23C41_GB20;
wire R27C1_GT10;
wire R24C24_GT10;
wire R26C20_GB40;
wire R13C28_GB50;
wire R15C45_GB50;
wire R14C35_GB70;
wire R28C16_W26;
wire R23C35_GB30;
wire R4C14_GB30;
wire R17C12_GB50;
wire R7C32_GB60;
wire R10C13_E81;
wire R4C30_GBO0;
wire R14C13_GB10;
wire R10C7_F5;
wire R28C13_W82;
wire R5C22_GB00;
wire R1C28_CE2;
wire R28C40_X06;
wire R22C6_GB50;
wire R1C47_N82;
wire R18C14_GB70;
wire R2C6_SPINE10;
wire R28C25_E11;
wire R17C32_GBO0;
wire R23C38_GB40;
wire R2C20_GB70;
wire R20C44_GBO1;
wire R10C43_W13;
wire R28C19_W11;
wire R22C11_GB50;
wire R11C44_GB00;
wire R15C22_GT00;
wire R13C32_GB00;
wire R22C45_GBO1;
wire R10C30_C5;
wire R16C3_GB30;
wire R1C32_E27;
wire R28C10_E10;
wire R18C15_GBO1;
wire R10C30_N27;
wire R9C11_GBO1;
wire R20C16_GB00;
wire R13C9_GT00;
wire R20C13_GB20;
wire R2C29_GT00;
wire R17C44_GB50;
wire R5C34_GT00;
wire R15C20_GB00;
wire R3C10_GB10;
wire R16C9_GB20;
wire R20C16_GB50;
wire R24C23_GB70;
wire R18C46_GBO0;
wire R5C36_GB30;
wire R28C16_X01;
wire R17C13_GT00;
wire R8C22_GB60;
wire R22C12_GB60;
wire R23C3_GB50;
wire R10C37_S80;
wire R28C40_D3;
wire R2C15_GB70;
wire R9C35_GB40;
wire R8C8_GB10;
wire R9C3_GT00;
wire R17C18_GB00;
wire R21C15_GT10;
wire R6C14_GB60;
wire R20C44_GB40;
wire R10C28_S80;
wire R28C34_W80;
wire R7C19_GB60;
wire R23C29_GB60;
wire R1C1_B3;
wire R10C37_LSR1;
wire R21C27_GB30;
wire R28C46_S23;
wire R20C19_SPINE21;
wire R17C27_GB30;
wire R26C45_GB10;
wire R10C37_Q6;
wire R21C24_GBO0;
wire R28C4_N20;
wire R28C43_A7;
wire R6C35_GB60;
wire R11C3_GB20;
wire R12C41_GB50;
wire R27C41_GB30;
wire R17C42_GBO1;
wire R11C14_GB60;
wire R10C27_S27;
wire R1C28_E25;
wire R13C39_GB50;
wire R2C45_GB50;
wire R10C16_Q7;
wire R20C33_GB10;
wire R28C10_F3;
wire R3C19_GBO0;
wire R17C25_GB30;
wire R14C11_GT00;
wire R26C28_GT10;
wire R21C20_GBO1;
wire R17C38_GT10;
wire R4C11_GBO0;
wire R8C19_GB50;
wire R27C7_GB60;
wire R15C12_GB60;
wire R13C45_GB20;
wire R1C1_LSR0;
wire R2C14_GB50;
wire R14C30_GB00;
wire R12C8_GB00;
wire R9C31_GT00;
wire R8C28_GB70;
wire R21C22_GB00;
wire R24C21_GB70;
wire R20C30_GT00;
wire R28C19_CLK0;
wire R28C43_Q2;
wire R8C6_GB50;
wire R9C5_GB00;
wire R2C16_GBO1;
wire R17C7_GB00;
wire R12C45_GB70;
wire R16C45_GB20;
wire R4C33_GB40;
wire R6C44_GT10;
wire R27C6_GB00;
wire R4C41_GB10;
wire R28C37_C3;
wire R28C34_E26;
wire R28C22_Q2;
wire R22C8_GB40;
wire R18C21_GB70;
wire R10C22_E12;
wire R6C26_GB10;
wire R17C9_GB70;
wire R28C19_B0;
wire R18C17_GBO0;
wire R7C17_GB00;
wire R5C2_GB40;
wire R4C41_GB50;
wire R17C38_GB60;
wire R10C30_S80;
wire R10C31_F6;
wire R9C37_GB30;
wire R25C9_GB20;
wire R7C14_GB20;
wire R8C34_GB30;
wire R21C41_GB50;
wire R10C19_SEL4;
wire R8C5_GB50;
wire R2C43_GB30;
wire R10C34_S25;
wire R15C15_GB00;
wire R5C41_GB50;
wire R25C11_GB70;
wire R10C19_W81;
wire R8C43_GB30;
wire R3C25_GT10;
wire R26C5_GB40;
wire R27C8_GB40;
wire R27C10_GB20;
wire R9C33_GB30;
wire R18C2_GB40;
wire R28C46_C0;
wire R14C42_GT00;
wire R22C15_GB50;
wire R4C17_GT00;
wire R26C24_GB70;
wire R10C31_S22;
wire R28C19_X01;
wire R12C27_GB40;
wire R24C20_GT00;
wire R7C17_GB10;
wire R17C18_GT00;
wire R13C4_GB30;
wire R13C17_GBO1;
wire R21C32_GB60;
wire R28C34_F0;
wire R28C43_E20;
wire R2C27_GB20;
wire R12C6_GB70;
wire R10C40_S20;
wire R21C40_GT00;
wire R25C21_GB50;
wire R13C16_GBO0;
wire R15C18_GB00;
wire R23C43_GB50;
wire R11C11_GB30;
wire R28C40_C2;
wire R12C43_GB70;
wire R1C47_X04;
wire R3C32_GB20;
wire R10C22_B4;
wire R10C13_N10;
wire R8C43_GT00;
wire R16C3_GB60;
wire R7C37_GB60;
wire R3C13_GB40;
wire R23C7_GBO1;
wire R10C37_SEL3;
wire R27C10_GBO0;
wire R11C6_GB60;
wire R27C16_GBO1;
wire R10C27_N83;
wire R10C29_S24;
wire R1C32_Q6;
wire R18C3_GB00;
wire R24C12_GB60;
wire R10C19_N10;
wire R2C19_GB00;
wire R14C5_GB00;
wire R24C41_GB30;
wire R3C46_GB70;
wire R5C42_GT00;
wire R27C7_GB10;
wire R26C34_GB70;
wire R8C32_GB30;
wire R23C19_GB40;
wire R28C40_S10;
wire R10C43_LSR0;
wire R10C19_S20;
wire R11C30_GBO0;
wire R14C17_GB50;
wire R10C27_E81;
wire R11C2_GB10;
wire R15C13_GB70;
wire R5C40_GB20;
wire R10C7_D2;
wire R28C34_C6;
wire R28C43_D0;
wire R17C29_GT10;
wire R9C24_GBO0;
wire R6C40_GB20;
wire R23C10_GB30;
wire R26C23_GB70;
wire R7C24_GT10;
wire R7C8_GB60;
wire R11C31_GB10;
wire R20C31_GB00;
wire R20C44_GB30;
wire R10C28_SEL2;
wire R27C11_GBO0;
wire R10C31_X05;
wire R20C9_GBO1;
wire R1C32_CE0;
wire R10C34_S24;
wire R28C22_W25;
wire R2C31_GB40;
wire R24C24_GB10;
wire R10C40_W27;
wire R28C19_S10;
wire R21C7_GBO0;
wire R27C13_GB20;
wire R28C43_S80;
wire R25C38_GB00;
wire R26C22_GB30;
wire R3C37_GB20;
wire R28C34_B0;
wire R6C24_GBO0;
wire R18C28_GB50;
wire R17C12_GB70;
wire R12C22_GB70;
wire R16C4_GT10;
wire R3C7_GB00;
wire R4C28_GB30;
wire R24C20_GB40;
wire R21C5_GB70;
wire R22C30_GBO1;
wire R29C28_Q7;
wire R11C33_GB20;
wire R8C13_GB30;
wire R1C32_F2;
wire R16C38_GBO1;
wire R1C32_W13;
wire R3C40_GB30;
wire R9C39_GT10;
wire R5C6_GT10;
wire R9C16_GB10;
wire R11C42_GB10;
wire R14C46_GBO0;
wire R10C25_W83;
wire R2C44_SPINE4;
wire R28C34_S83;
wire R2C24_GB00;
wire R8C34_GB60;
wire R11C15_GB70;
wire R3C39_GB30;
wire R9C13_GB00;
wire R23C24_GBO0;
wire R3C8_GB40;
wire R20C5_GT10;
wire R12C24_GB20;
wire R10C31_W83;
wire R14C6_GB30;
wire R10C22_CLK2;
wire R4C38_GB40;
wire R22C28_GT10;
wire R15C40_GB40;
wire R21C44_GB70;
wire R18C21_GB30;
wire R25C12_GB20;
wire R1C47_SN20;
wire R2C37_GBO1;
wire R22C30_GT00;
wire R23C2_GB50;
wire R22C33_GB00;
wire R1C32_W23;
wire R10C19_W83;
wire R10C43_Q6;
wire R15C43_GBO1;
wire R18C10_GB00;
wire R15C14_GB20;
wire R21C8_GB70;
wire R2C30_GB40;
wire R28C37_B6;
wire R4C18_GB10;
wire R1C28_N81;
wire R10C22_SEL1;
wire R27C34_GB20;
wire R3C32_GB00;
wire R18C24_GB70;
wire R21C32_GB40;
wire R17C12_GB00;
wire R11C24_GB40;
wire R17C22_GBO1;
wire R1C47_SEL7;
wire R17C9_GT10;
wire R6C23_GB60;
wire R2C35_GBO1;
wire R28C34_SN20;
wire R18C43_GT10;
wire R9C41_GB70;
wire R10C30_SEL7;
wire R8C28_GB40;
wire R18C19_GT10;
wire R29C28_LSR0;
wire R13C17_GT00;
wire R5C20_GB20;
wire R10C34_E20;
wire R28C19_SEL3;
wire R10C37_W12;
wire R2C46_GT00;
wire R20C25_GBO0;
wire R24C3_GB70;
wire R28C46_S12;
wire R21C13_GBO0;
wire R2C29_GB70;
wire R7C25_GB20;
wire R14C22_GB40;
wire R12C6_GT00;
wire R2C26_GB70;
wire R15C17_GB60;
wire R10C34_CLK1;
wire R15C35_GB20;
wire R1C32_SEL3;
wire R1C47_CLK0;
wire R9C44_GB10;
wire R1C47_Q1;
wire R2C32_GB60;
wire R22C35_GB40;
wire R24C45_GB30;
wire R2C23_SPINE9;
wire R3C39_GT00;
wire R18C15_GBO0;
wire R6C26_GB20;
wire R21C37_GT10;
wire R3C4_GBO0;
wire R20C25_GT00;
wire R22C27_GT10;
wire R5C25_GB30;
wire R27C32_GB10;
wire R20C32_SPINE24;
wire R10C10_S81;
wire R28C13_F1;
wire R27C41_GT10;
wire R9C20_GB00;
wire R18C40_GT00;
wire R7C14_GB50;
wire R12C3_GB70;
wire R28C43_SEL1;
wire R26C34_GBO0;
wire R23C45_GT00;
wire R6C19_GB10;
wire R25C45_GBO0;
wire R15C30_GT10;
wire R12C34_GB20;
wire R26C11_GB50;
wire R26C17_GBO1;
wire R11C38_GB20;
wire R15C39_GB40;
wire R1C32_E22;
wire R10C37_C6;
wire R10C10_X03;
wire R28C31_SEL6;
wire R14C4_GB20;
wire R28C43_D7;
wire R22C27_GT00;
wire R10C10_EW20;
wire R10C22_Q6;
wire R13C43_GT10;
wire R10C29_E11;
wire R5C19_GT10;
wire R20C15_GB60;
wire R27C39_GB40;
wire R7C8_GT10;
wire R2C22_GB60;
wire R10C22_Q4;
wire R3C15_GB30;
wire R11C26_GB60;
wire R2C23_GB40;
wire R6C5_GT10;
wire R10C28_N25;
wire R15C8_GB40;
wire R10C13_E80;
wire R27C20_GB50;
wire R28C19_N22;
wire R2C31_GB10;
wire R15C19_GB10;
wire R10C25_EW10;
wire R28C10_N10;
wire R4C17_GB10;
wire R26C44_GB50;
wire R4C31_GBO1;
wire R26C43_GBO1;
wire R10C43_N10;
wire R25C13_GBO0;
wire R28C28_Q7;
wire R5C2_GB60;
wire R2C17_GT10;
wire R14C28_GB70;
wire R9C45_GB60;
wire R23C36_GBO0;
wire R6C13_GBO1;
wire R10C29_X03;
wire R12C21_GB40;
wire R28C28_W80;
wire R28C40_E83;
wire R28C13_Q2;
wire R25C37_GB00;
wire R15C22_GB40;
wire R20C4_GB10;
wire R3C5_GB30;
wire R12C1_GBO0;
wire R7C39_GB70;
wire R23C45_GB40;
wire R1C28_C1;
wire R10C19_X08;
wire R14C17_GB30;
wire R1C32_SEL1;
wire R28C28_SEL6;
wire R28C10_E23;
wire R21C21_GT00;
wire R23C4_GB60;
wire R10C13_S21;
wire R1C47_Q5;
wire R28C31_F6;
wire R22C21_GBO1;
wire R23C12_GB40;
wire R9C25_GB60;
wire R2C24_GB70;
wire R16C45_GB30;
wire R28C22_D4;
wire R12C38_GB10;
wire R28C25_Q4;
wire R10C22_Q3;
wire R28C43_A1;
wire R21C28_GB70;
wire R3C9_GB00;
wire R14C2_GB40;
wire R3C24_GT00;
wire R17C24_GT10;
wire R4C5_GBO0;
wire R10C25_Q4;
wire R21C20_GT00;
wire R11C9_GB20;
wire R28C16_B7;
wire R16C30_GBO0;
wire R22C4_GB50;
wire R16C16_GB70;
wire R5C28_GT00;
wire R6C28_GT10;
wire R25C6_GT10;
wire R6C21_GB70;
wire R26C7_GBO1;
wire R2C15_SPINE13;
wire R7C27_GB50;
wire R16C16_GBO0;
wire R7C36_GB40;
wire R27C46_GB00;
wire R26C40_GB40;
wire R5C1_GBO1;
wire R9C30_GB00;
wire R26C18_GB30;
wire R10C25_Q2;
wire R25C1_GT00;
wire R6C37_GB70;
wire R15C30_GB50;
wire R28C10_S25;
wire R26C45_GT10;
wire R10C31_E23;
wire R25C26_GB10;
wire R11C41_GB50;
wire R7C9_GB50;
wire R5C15_GB30;
wire R16C8_GB50;
wire R4C40_GBO0;
wire R9C35_GB50;
wire R10C7_X06;
wire R9C19_GB20;
wire R24C40_GB10;
wire R20C12_GB40;
wire R3C42_GB00;
wire R9C13_GT00;
wire R4C7_GT00;
wire R7C15_GT10;
wire R16C28_GT10;
wire R3C46_GT10;
wire R6C6_GB50;
wire R10C30_W10;
wire R10C26_W11;
wire R22C2_GB00;
wire R1C32_F7;
wire R3C43_GBO1;
wire R1C47_EW10;
wire R4C34_GB50;
wire R2C31_GB60;
wire R23C39_GT10;
wire R10C16_A4;
wire R9C17_GB00;
wire R23C37_GB10;
wire R2C37_GT10;
wire R12C2_GB50;
wire R28C25_A3;
wire R2C39_SPINE5;
wire R23C24_GT00;
wire R27C25_GB10;
wire R17C35_GB40;
wire R27C20_GT00;
wire R14C38_GB50;
wire R10C26_N80;
wire R15C9_GB70;
wire R12C28_GB50;
wire R10C40_E24;
wire R4C15_GBO0;
wire R7C8_GB00;
wire R16C25_GB40;
wire R11C26_GBO1;
wire R20C13_GB70;
wire R26C19_GB00;
wire R10C40_C0;
wire R22C2_GT10;
wire R7C42_GB70;
wire R5C18_GB30;
wire R20C27_GB30;
wire R5C9_GB70;
wire R12C29_GB70;
wire R1C1_W82;
wire R17C19_GBO1;
wire R1C1_X06;
wire R26C21_GBO0;
wire R23C2_GT00;
wire R8C19_GBO0;
wire R10C30_E81;
wire R27C23_GB00;
wire R3C19_GB10;
wire R26C2_GB40;
wire R6C37_GB50;
wire R21C34_GB30;
wire R9C23_GB60;
wire R20C14_GBO0;
wire R16C23_GB40;
wire R13C33_GBO1;
wire R10C7_B7;
wire R25C31_GT00;
wire R28C10_N83;
wire R24C26_GB20;
wire R5C32_GB40;
wire R25C5_GB50;
wire R2C21_GT10;
wire R10C34_S10;
wire R14C38_GT00;
wire R14C33_GB60;
wire R12C14_GB60;
wire R7C31_GB20;
wire R13C26_GT10;
wire R20C8_GB10;
wire R20C35_GT10;
wire R23C36_GB30;
wire R14C5_GT10;
wire R10C22_E11;
wire R28C4_N21;
wire R23C25_GB40;
wire R10C13_S81;
wire R9C14_GBO1;
wire R23C23_GB00;
wire R13C42_GBO0;
wire R20C27_GT10;
wire R4C15_GB30;
wire R17C33_GBO0;
wire R2C22_GT00;
wire R17C22_GB60;
wire R23C3_GBO1;
wire R28C28_C5;
wire R15C40_GB20;
wire R1C28_E21;
wire R28C31_SEL3;
wire R23C40_GB00;
wire R14C43_GB00;
wire R20C30_GB30;
wire R13C5_GT10;
wire R10C13_F4;
wire R28C40_S27;
wire R26C8_GB10;
wire R20C42_GB00;
wire R8C18_GB00;
wire R9C31_GB60;
wire R11C8_GT00;
wire R11C13_GB20;
wire R27C28_GB70;
wire R27C16_GT00;
wire R9C33_GB20;
wire R10C34_S13;
wire R25C43_GB10;
wire R8C11_GT00;
wire R11C2_GB00;
wire R17C41_GBO0;
wire R10C37_A1;
wire R22C40_GT10;
wire R13C30_GT00;
wire R10C40_D1;
wire R28C7_W21;
wire R23C2_GT10;
wire R23C31_GT10;
wire R10C25_W22;
wire R28C10_B0;
wire R3C14_GB50;
wire R6C27_GB00;
wire R2C1_GBO0;
wire R26C34_GB50;
wire R1C47_E11;
wire R28C46_Q7;
wire R27C35_GT00;
wire R10C27_S25;
wire R28C37_W10;
wire R29C28_N27;
wire R24C7_GB40;
wire R10C30_C2;
wire R8C12_GBO0;
wire R21C15_GB30;
wire R9C42_GB50;
wire R6C5_GB40;
wire R15C12_GB40;
wire R4C43_GB00;
wire R10C26_F3;
wire R6C13_GB70;
wire R15C11_GT00;
wire R14C27_GB00;
wire R22C33_GB30;
wire R23C2_GB20;
wire R11C28_GB40;
wire R28C43_A5;
wire R17C17_GB70;
wire R16C36_GBO1;
wire R15C30_GB70;
wire R21C8_GB60;
wire R6C6_GT00;
wire R2C35_SPINE1;
wire R20C20_GB40;
wire R25C24_GT00;
wire R6C2_GB10;
wire R2C16_GB30;
wire R25C39_GT10;
wire R3C26_GB50;
wire R24C3_GB20;
wire R24C32_GBO1;
wire R10C40_A2;
wire R3C46_GB20;
wire R1C1_LSR2;
wire R5C14_GB40;
wire R6C45_GB10;
wire R13C25_GBO0;
wire R6C12_GB50;
wire R23C43_GBO0;
wire R28C37_S21;
wire R9C38_GB00;
wire R20C23_GT00;
wire R25C42_GT00;
wire R17C8_GBO1;
wire R2C10_GB50;
wire R13C20_GB00;
wire R21C24_GB20;
wire R28C22_X02;
wire R10C37_W24;
wire R15C16_GB00;
wire R26C22_GB50;
wire R28C25_SEL3;
wire R7C33_GB50;
wire R13C43_GB00;
wire R27C20_GB70;
wire R18C41_GT10;
wire R10C40_B4;
wire R13C31_GB10;
wire R24C37_GB60;
wire R10C19_CLK0;
wire R28C28_W22;
wire R6C41_GB70;
wire R11C37_GT00;
wire R20C29_GB40;
wire R13C12_GB70;
wire R10C30_UNK122;
wire R5C31_GT00;
wire R9C32_GT00;
wire R22C16_GB20;
wire R17C25_GB70;
wire R23C32_GBO0;
wire R10C7_W13;
wire R10C7_E11;
wire R10C43_S24;
wire R28C13_B4;
wire R28C13_D0;
wire R16C21_GT00;
wire R28C40_Q3;
wire R2C13_GB10;
wire R10C27_S82;
wire R20C4_SPINE16;
wire R27C13_GT00;
wire R20C10_GT00;
wire R3C14_GB20;
wire R28C10_W10;
wire R22C28_GB70;
wire R28C13_X08;
wire R18C5_GT00;
wire R23C29_GB30;
wire R17C31_GB50;
wire R10C26_Q4;
wire R2C8_GB00;
wire R28C7_SEL6;
wire R24C29_GT00;
wire R10C31_D7;
wire R3C7_GB40;
wire R22C37_GB10;
wire R18C5_GBO0;
wire R28C43_B4;
wire R10C27_CE0;
wire R28C28_S13;
wire R11C41_GBO0;
wire R2C42_GBO1;
wire R20C46_GT00;
wire R27C32_GBO0;
wire R18C10_GB50;
wire R17C18_GB20;
wire R28C25_C0;
wire R5C26_GB40;
wire R16C1_GT00;
wire R4C27_GB50;
wire R4C23_GB20;
wire R7C9_GB40;
wire R2C2_GB70;
wire R27C41_GB60;
wire R13C37_GBO1;
wire R28C13_E27;
wire R2C24_SPINE12;
wire R1C47_Q2;
wire R20C3_GB10;
wire R27C2_GB50;
wire R13C22_GB50;
wire R25C24_GT10;
wire R1C28_N27;
wire R10C19_W13;
wire R28C34_W21;
wire R9C6_GB70;
wire R8C17_GB00;
wire R10C43_S12;
wire R25C8_GB20;
wire R26C34_GB30;
wire R21C4_GB00;
wire R16C42_GB30;
wire R20C14_GT10;
wire R2C20_GT10;
wire R1C28_S25;
wire R14C37_GBO0;
wire R25C46_GB50;
wire R18C1_GBO1;
wire R5C37_GB10;
wire R11C17_GB30;
wire R10C29_D5;
wire R13C43_GB50;
wire R14C21_GB10;
wire R16C28_GB40;
wire R9C37_GB50;
wire R22C22_GB50;
wire R23C46_GB60;
wire R27C44_GB10;
wire R10C29_C1;
wire R28C7_N11;
wire R10C28_CLK2;
wire R10C7_CE0;
wire R23C46_GT00;
wire R9C29_GB30;
wire R23C44_GB20;
wire R2C20_GB50;
wire R10C28_S27;
wire R10C31_S25;
wire R10C37_W13;
wire R10C28_Q7;
wire R21C21_GB00;
wire R9C14_GB50;
wire R25C8_GB30;
wire R7C2_GT00;
wire R16C40_GBO0;
wire R10C34_S22;
wire R10C37_B6;
wire R28C19_E20;
wire R21C43_GB30;
wire R3C26_GB70;
wire R4C36_GB20;
wire R26C41_GB00;
wire R2C21_GB70;
wire R15C34_GBO0;
wire R7C38_GB60;
wire R17C21_GT10;
wire R16C1_GT10;
wire R18C26_GT10;
wire R15C6_GB20;
wire R24C43_GB50;
wire R14C5_GBO1;
wire R1C1_S27;
wire R2C10_SPINE10;
wire R23C12_GB70;
wire R12C37_GT10;
wire R8C28_GB20;
wire R10C27_W82;
wire R5C7_GBO0;
wire R11C25_GB40;
wire R10C28_SPINE17;
wire R18C44_GT10;
wire R17C19_GB10;
wire R22C42_GB40;
wire R10C26_W25;
wire R12C16_GB60;
wire R28C46_W22;
wire R28C31_CLK1;
wire R18C20_GB60;
wire R3C42_GT00;
wire R10C30_UNK125;
wire R12C36_GB20;
wire R17C35_GT00;
wire R1C1_SEL6;
wire R14C36_GB00;
wire R20C44_GT10;
wire R28C31_Q5;
wire R7C21_GB70;
wire R20C15_GB40;
wire R1C47_LSR0;
wire R20C37_GT10;
wire R9C43_GB50;
wire R4C23_GB10;
wire R4C46_GB40;
wire R22C7_GB10;
wire R15C46_GBO1;
wire R10C29_N83;
wire R5C12_GBO0;
wire R10C40_N24;
wire R28C7_SEL3;
wire R10C40_D2;
wire R14C34_GB20;
wire R28C31_F0;
wire R29C28_N21;
wire R26C14_GB40;
wire R16C25_GB70;
wire R3C22_GT00;
wire R26C21_GT10;
wire R3C5_GB10;
wire R10C30_S27;
wire R10C37_W10;
wire R18C13_GB60;
wire R28C46_S13;
wire R23C9_GB60;
wire R11C18_GT00;
wire R10C30_D3;
wire R15C24_GB30;
wire R13C13_GB70;
wire R26C15_GT10;
wire R10C28_S26;
wire R16C31_GB20;
wire R3C2_GB00;
wire R12C8_GBO1;
wire R28C13_E83;
wire R3C17_GB60;
wire R3C1_GBO1;
wire R10C40_LSR0;
wire R11C27_GB40;
wire R7C2_GBO0;
wire R16C18_GB20;
wire R22C22_GB40;
wire R28C22_EW20;
wire R1C47_B7;
wire R10C16_D2;
wire R28C43_SN20;
wire R7C17_GB40;
wire R28C13_Q4;
wire R28C22_SN10;
wire R10C22_C7;
wire R17C4_GB10;
wire R10C7_N12;
wire R5C19_GB00;
wire R23C17_GB00;
wire R21C20_GB20;
wire R28C19_B5;
wire R5C34_GB40;
wire R12C17_GB30;
wire R10C22_S82;
wire R28C19_S21;
wire R3C32_GT00;
wire R4C41_GBO0;
wire R10C13_F6;
wire R16C5_GB30;
wire R10C27_E23;
wire R18C7_GB60;
wire R1C1_B6;
wire R1C1_N12;
wire R10C30_SEL6;
wire R9C12_GB20;
wire R22C28_GB50;
wire R28C43_B7;
wire R28C4_A0;
wire R2C33_GBO1;
wire R10C27_E27;
wire R7C17_GB60;
wire R18C41_GBO0;
wire R10C34_X06;
wire R22C31_GT10;
wire R15C2_GB10;
wire R18C4_GB20;
wire R21C4_GBO1;
wire R26C33_GB50;
wire R21C17_GB10;
wire R14C23_GBO0;
wire R23C4_GBO1;
wire R18C24_GBO0;
wire R15C43_GB10;
wire R1C47_F4;
wire R5C17_GBO1;
wire R3C21_GBO1;
wire R13C25_GB40;
wire R13C28_GT10;
wire R26C37_GB10;
wire R28C37_E22;
wire R14C26_GB20;
wire R18C39_GB00;
wire R26C42_GB60;
wire R9C38_GB10;
wire R10C25_N23;
wire R2C26_GB00;
wire R28C37_D1;
wire R5C21_GB50;
wire R17C42_GB40;
wire R3C22_GB10;
wire R13C13_GT00;
wire R28C10_E20;
wire R25C16_GB70;
wire R17C45_GB00;
wire R17C15_GB70;
wire R4C46_GBO0;
wire R9C41_GB30;
wire R11C43_GT10;
wire R20C42_GT00;
wire R15C35_GB10;
wire R20C23_GB70;
wire R25C38_GB60;
wire R17C27_GB60;
wire R28C16_S20;
wire R11C43_GBO0;
wire R6C18_GB50;
wire R13C6_GB10;
wire R4C27_GT10;
wire R20C46_GB60;
wire R16C36_GBO0;
wire R21C31_GBO1;
wire R25C18_GB40;
wire R2C16_GT00;
wire R15C14_GT00;
wire R1C32_E20;
wire R14C37_GB10;
wire R24C37_GT10;
wire R21C17_GBO0;
wire R23C29_GB70;
wire R4C26_GBO0;
wire R10C25_A3;
wire R7C8_GB40;
wire R3C11_GB70;
wire R10C19_N83;
wire R28C10_E12;
wire R26C40_GB30;
wire R10C7_S25;
wire R20C27_GB60;
wire R28C10_E83;
wire R28C37_N80;
wire R18C46_GB30;
wire R24C31_GB00;
wire R10C13_S12;
wire R10C26_A7;
wire R24C45_GB40;
wire R16C12_GB40;
wire R4C5_GBO1;
wire R16C38_GB00;
wire R20C30_GBO1;
wire R1C1_C7;
wire R17C42_GB10;
wire R5C34_GB00;
wire R10C16_S26;
wire R16C34_GT00;
wire R13C8_GB00;
wire R10C28_W12;
wire R5C28_GT10;
wire R12C16_GB00;
wire R11C33_GT00;
wire R24C34_GB70;
wire R26C28_GB30;
wire R4C38_GBO1;
wire R16C29_GB30;
wire R17C30_GB30;
wire R17C26_GT00;
wire R10C22_SN20;
wire R10C31_N23;
wire R28C4_N82;
wire R3C40_GB20;
wire R14C5_GB40;
wire R23C21_GB50;
wire R13C14_GB20;
wire R21C15_GB60;
wire R20C39_GT10;
wire R23C20_GBO0;
wire R13C36_GBO1;
wire R10C13_N20;
wire R11C24_GB60;
wire R5C42_GB70;
wire R23C42_GB10;
wire R10C10_SEL3;
wire R28C40_SEL1;
wire R27C5_GB10;
wire R11C22_GB10;
wire R9C15_GB00;
wire R10C22_F7;
wire R23C5_GT00;
wire R21C15_GB50;
wire R10C13_X08;
wire R13C9_GB20;
wire R15C27_GB50;
wire R1C47_B6;
wire R13C15_GBO1;
wire R10C43_A1;
wire R1C32_S24;
wire R25C21_GB70;
wire R15C43_GB50;
wire R26C40_GB50;
wire R17C15_GBO1;
wire R3C13_GBO1;
wire R16C42_GB60;
wire R18C15_GT00;
wire R10C19_SEL1;
wire R2C33_SPINE3;
wire R20C24_GB50;
wire R20C8_GBO0;
wire R28C22_D2;
wire R28C43_S10;
wire R14C20_GT00;
wire R18C3_GB50;
wire R16C42_GT00;
wire R17C22_GB70;
wire R24C22_GBO1;
wire R16C43_GB70;
wire R2C33_GB70;
wire R6C17_GB00;
wire R5C4_GBO1;
wire R2C18_GB40;
wire R23C16_GBO0;
wire R4C32_GB30;
wire R3C41_GBO1;
wire R28C34_S81;
wire R10C16_Q4;
wire R15C32_GT00;
wire R24C23_GB20;
wire R22C19_GT10;
wire R27C43_GB10;
wire R8C19_GT10;
wire R10C34_B2;
wire R10C37_N80;
wire R27C9_GB40;
wire R3C35_GBO0;
wire R28C10_S21;
wire R6C8_GB00;
wire R28C31_N26;
wire R28C37_C0;
wire R7C25_GB00;
wire R2C35_GT10;
wire R28C28_W20;
wire R16C6_GB00;
wire R12C21_GT00;
wire R21C26_GB50;
wire R8C35_GB70;
wire R11C27_GB50;
wire R28C40_CLK1;
wire R24C29_GT10;
wire R9C32_GB20;
wire R20C29_GBO0;
wire R10C22_X07;
wire R10C28_N24;
wire R27C4_GB30;
wire R24C38_GB00;
wire R20C18_GB60;
wire R21C37_GB20;
wire R27C42_GB40;
wire R10C25_W25;
wire R5C18_GT00;
wire R27C8_GB60;
wire R10C30_X04;
wire R8C14_GB00;
wire R25C29_GB10;
wire R28C43_CE2;
wire R9C24_GBO1;
wire R28C34_X02;
wire R7C15_GB40;
wire R28C31_S12;
wire R12C43_GB00;
wire R7C9_GB00;
wire R28C34_S13;
wire R1C1_F1;
wire R16C10_GB10;
wire R4C13_GB10;
wire R28C13_W12;
wire R6C36_GT10;
wire R17C22_GB30;
wire R25C29_GBO0;
wire R11C45_GB30;
wire R14C8_GB20;
wire R23C25_GB60;
wire R10C29_SEL0;
wire R28C4_F5;
wire R28C13_N81;
wire R28C25_Q5;
wire R22C13_GB30;
wire R24C37_GBO1;
wire R1C32_F4;
wire R27C20_GB00;
wire R17C8_GB10;
wire R5C32_GB50;
wire R1C47_D3;
wire R8C30_GB10;
wire R7C41_GB30;
wire R2C31_GB30;
wire R26C2_GB00;
wire R10C16_W10;
wire R25C7_GB70;
wire R28C4_B1;
wire R28C37_S23;
wire R28C7_X04;
wire R25C44_GB50;
wire R24C20_GB10;
wire R10C7_F1;
wire R14C17_GT00;
wire R13C16_GB70;
wire R22C13_GB10;
wire R21C28_GB60;
wire R21C36_GB60;
wire R17C20_GB20;
wire R27C27_GB50;
wire R6C5_GBO1;
wire R6C41_GBO0;
wire R8C30_GB40;
wire R29C28_N82;
wire R22C23_GB20;
wire R23C11_GB20;
wire R4C23_GB30;
wire R10C29_S26;
wire R23C40_GT10;
wire R2C8_GB10;
wire R25C10_GB70;
wire R6C31_GB00;
wire R10C40_S11;
wire R29C28_Q4;
wire R10C29_C7;
wire R10C40_W11;
wire R12C46_GB30;
wire R3C44_GB70;
wire R12C42_GB10;
wire R10C43_F3;
wire R3C20_GB30;
wire R1C28_SN20;
wire R27C25_GBO0;
wire R2C28_GB60;
wire R1C47_N81;
wire R7C28_GT00;
wire R10C31_B1;
wire R9C25_GT10;
wire R17C25_GB00;
wire R20C29_GB50;
wire R25C12_GB40;
wire R4C43_GB20;
wire R7C45_GB30;
wire R13C30_GBO1;
wire R28C10_F2;
wire R18C45_GT10;
wire R3C12_GT00;
wire R5C19_GBO1;
wire R17C16_GBO0;
wire R1C32_D5;
wire R10C22_CLK0;
wire R28C16_S21;
wire R17C42_GT00;
wire R4C17_GB40;
wire R1C1_S26;
wire R6C24_GB20;
assign R10C27_UNK127 = R9C47_F6;
assign R10C27_UNK124 = R29C29_F6;
assign R10C27_UNK126 = R15C1_F6;
assign R10C27_UNK125 = R9C1_F6;
assign R10C27_UNK128 = R17C47_F6;
assign R10C27_UNK123 = R29C28_F6;
assign R10C27_UNK121 = R1C28_F6;
assign R10C27_UNK122 = R1C29_F6;
assign R10C28_UNK127 = R9C47_F6;
assign R10C28_UNK124 = R29C29_F6;
assign R10C28_UNK126 = R15C1_F6;
assign R10C28_UNK125 = R9C1_F6;
assign R10C28_UNK128 = R17C47_F6;
assign R10C28_UNK123 = R29C28_F6;
assign R10C28_UNK121 = R1C28_F6;
assign R10C28_UNK122 = R1C29_F6;
assign R10C30_UNK127 = R9C47_F6;
assign R10C30_UNK124 = R29C29_F6;
assign R10C30_UNK126 = R15C1_F6;
assign R10C30_UNK125 = R9C1_F6;
assign R10C30_UNK128 = R17C47_F6;
assign R10C30_UNK123 = R29C28_F6;
assign R10C30_UNK121 = R1C28_F6;
assign R10C30_UNK122 = R1C29_F6;
assign R10C29_UNK127 = R9C47_F6;
assign R10C29_UNK124 = R29C29_F6;
assign R10C29_UNK126 = R15C1_F6;
assign R10C29_UNK125 = R9C1_F6;
assign R10C29_UNK128 = R17C47_F6;
assign R10C29_UNK123 = R29C28_F6;
assign R10C29_UNK121 = R1C28_F6;
assign R10C29_UNK122 = R1C29_F6;
assign R2C4_SPINE8 = R10C27_SPINE8;
assign R2C8_SPINE8 = R10C27_SPINE8;
assign R2C12_SPINE8 = R10C27_SPINE8;
assign R2C16_SPINE8 = R10C27_SPINE8;
assign R2C20_SPINE8 = R10C27_SPINE8;
assign R2C24_SPINE8 = R10C27_SPINE8;
assign R2C3_SPINE9 = R10C27_SPINE9;
assign R2C7_SPINE9 = R10C27_SPINE9;
assign R2C11_SPINE9 = R10C27_SPINE9;
assign R2C15_SPINE9 = R10C27_SPINE9;
assign R2C19_SPINE9 = R10C27_SPINE9;
assign R2C23_SPINE9 = R10C27_SPINE9;
assign R2C27_SPINE9 = R10C27_SPINE9;
assign R2C2_SPINE10 = R10C27_SPINE10;
assign R2C6_SPINE10 = R10C27_SPINE10;
assign R2C10_SPINE10 = R10C27_SPINE10;
assign R2C14_SPINE10 = R10C27_SPINE10;
assign R2C18_SPINE10 = R10C27_SPINE10;
assign R2C22_SPINE10 = R10C27_SPINE10;
assign R2C26_SPINE10 = R10C27_SPINE10;
assign R2C1_SPINE11 = R10C27_SPINE11;
assign R2C5_SPINE11 = R10C27_SPINE11;
assign R2C9_SPINE11 = R10C27_SPINE11;
assign R2C13_SPINE11 = R10C27_SPINE11;
assign R2C17_SPINE11 = R10C27_SPINE11;
assign R2C21_SPINE11 = R10C27_SPINE11;
assign R2C25_SPINE11 = R10C27_SPINE11;
assign R2C4_SPINE12 = R10C27_SPINE12;
assign R2C8_SPINE12 = R10C27_SPINE12;
assign R2C12_SPINE12 = R10C27_SPINE12;
assign R2C16_SPINE12 = R10C27_SPINE12;
assign R2C20_SPINE12 = R10C27_SPINE12;
assign R2C24_SPINE12 = R10C27_SPINE12;
assign R2C3_SPINE13 = R10C27_SPINE13;
assign R2C7_SPINE13 = R10C27_SPINE13;
assign R2C11_SPINE13 = R10C27_SPINE13;
assign R2C15_SPINE13 = R10C27_SPINE13;
assign R2C19_SPINE13 = R10C27_SPINE13;
assign R2C23_SPINE13 = R10C27_SPINE13;
assign R2C27_SPINE13 = R10C27_SPINE13;
assign R20C4_SPINE16 = R10C28_SPINE16;
assign R20C8_SPINE16 = R10C28_SPINE16;
assign R20C12_SPINE16 = R10C28_SPINE16;
assign R20C16_SPINE16 = R10C28_SPINE16;
assign R20C20_SPINE16 = R10C28_SPINE16;
assign R20C24_SPINE16 = R10C28_SPINE16;
assign R20C3_SPINE17 = R10C28_SPINE17;
assign R20C7_SPINE17 = R10C28_SPINE17;
assign R20C11_SPINE17 = R10C28_SPINE17;
assign R20C15_SPINE17 = R10C28_SPINE17;
assign R20C19_SPINE17 = R10C28_SPINE17;
assign R20C23_SPINE17 = R10C28_SPINE17;
assign R20C27_SPINE17 = R10C28_SPINE17;
assign R20C2_SPINE18 = R10C28_SPINE18;
assign R20C6_SPINE18 = R10C28_SPINE18;
assign R20C10_SPINE18 = R10C28_SPINE18;
assign R20C14_SPINE18 = R10C28_SPINE18;
assign R20C18_SPINE18 = R10C28_SPINE18;
assign R20C22_SPINE18 = R10C28_SPINE18;
assign R20C26_SPINE18 = R10C28_SPINE18;
assign R20C1_SPINE19 = R10C28_SPINE19;
assign R20C5_SPINE19 = R10C28_SPINE19;
assign R20C9_SPINE19 = R10C28_SPINE19;
assign R20C13_SPINE19 = R10C28_SPINE19;
assign R20C17_SPINE19 = R10C28_SPINE19;
assign R20C21_SPINE19 = R10C28_SPINE19;
assign R20C25_SPINE19 = R10C28_SPINE19;
assign R20C4_SPINE20 = R10C28_SPINE20;
assign R20C8_SPINE20 = R10C28_SPINE20;
assign R20C12_SPINE20 = R10C28_SPINE20;
assign R20C16_SPINE20 = R10C28_SPINE20;
assign R20C20_SPINE20 = R10C28_SPINE20;
assign R20C24_SPINE20 = R10C28_SPINE20;
assign R20C3_SPINE21 = R10C28_SPINE21;
assign R20C7_SPINE21 = R10C28_SPINE21;
assign R20C11_SPINE21 = R10C28_SPINE21;
assign R20C15_SPINE21 = R10C28_SPINE21;
assign R20C19_SPINE21 = R10C28_SPINE21;
assign R20C23_SPINE21 = R10C28_SPINE21;
assign R20C27_SPINE21 = R10C28_SPINE21;
assign R2C32_SPINE0 = R10C30_SPINE0;
assign R2C36_SPINE0 = R10C30_SPINE0;
assign R2C40_SPINE0 = R10C30_SPINE0;
assign R2C44_SPINE0 = R10C30_SPINE0;
assign R2C31_SPINE1 = R10C30_SPINE1;
assign R2C35_SPINE1 = R10C30_SPINE1;
assign R2C39_SPINE1 = R10C30_SPINE1;
assign R2C43_SPINE1 = R10C30_SPINE1;
assign R2C30_SPINE2 = R10C30_SPINE2;
assign R2C34_SPINE2 = R10C30_SPINE2;
assign R2C38_SPINE2 = R10C30_SPINE2;
assign R2C42_SPINE2 = R10C30_SPINE2;
assign R2C46_SPINE2 = R10C30_SPINE2;
assign R2C29_SPINE3 = R10C30_SPINE3;
assign R2C33_SPINE3 = R10C30_SPINE3;
assign R2C37_SPINE3 = R10C30_SPINE3;
assign R2C41_SPINE3 = R10C30_SPINE3;
assign R2C45_SPINE3 = R10C30_SPINE3;
assign R2C32_SPINE4 = R10C30_SPINE4;
assign R2C36_SPINE4 = R10C30_SPINE4;
assign R2C40_SPINE4 = R10C30_SPINE4;
assign R2C44_SPINE4 = R10C30_SPINE4;
assign R2C31_SPINE5 = R10C30_SPINE5;
assign R2C35_SPINE5 = R10C30_SPINE5;
assign R2C39_SPINE5 = R10C30_SPINE5;
assign R2C43_SPINE5 = R10C30_SPINE5;
assign R20C32_SPINE24 = R10C29_SPINE24;
assign R20C36_SPINE24 = R10C29_SPINE24;
assign R20C40_SPINE24 = R10C29_SPINE24;
assign R20C44_SPINE24 = R10C29_SPINE24;
assign R20C31_SPINE25 = R10C29_SPINE25;
assign R20C35_SPINE25 = R10C29_SPINE25;
assign R20C39_SPINE25 = R10C29_SPINE25;
assign R20C43_SPINE25 = R10C29_SPINE25;
assign R20C30_SPINE26 = R10C29_SPINE26;
assign R20C34_SPINE26 = R10C29_SPINE26;
assign R20C38_SPINE26 = R10C29_SPINE26;
assign R20C42_SPINE26 = R10C29_SPINE26;
assign R20C46_SPINE26 = R10C29_SPINE26;
assign R20C29_SPINE27 = R10C29_SPINE27;
assign R20C33_SPINE27 = R10C29_SPINE27;
assign R20C37_SPINE27 = R10C29_SPINE27;
assign R20C41_SPINE27 = R10C29_SPINE27;
assign R20C45_SPINE27 = R10C29_SPINE27;
assign R20C32_SPINE28 = R10C29_SPINE28;
assign R20C36_SPINE28 = R10C29_SPINE28;
assign R20C40_SPINE28 = R10C29_SPINE28;
assign R20C44_SPINE28 = R10C29_SPINE28;
assign R20C31_SPINE29 = R10C29_SPINE29;
assign R20C35_SPINE29 = R10C29_SPINE29;
assign R20C39_SPINE29 = R10C29_SPINE29;
assign R20C43_SPINE29 = R10C29_SPINE29;
assign R3C1_GT00 = R2C1_GT00;
assign R3C1_GT10 = R2C1_GT10;
assign R4C1_GT00 = R2C1_GT00;
assign R4C1_GT10 = R2C1_GT10;
assign R5C1_GT00 = R2C1_GT00;
assign R5C1_GT10 = R2C1_GT10;
assign R6C1_GT00 = R2C1_GT00;
assign R6C1_GT10 = R2C1_GT10;
assign R7C1_GT00 = R2C1_GT00;
assign R7C1_GT10 = R2C1_GT10;
assign R8C1_GT00 = R2C1_GT00;
assign R8C1_GT10 = R2C1_GT10;
assign R9C1_GT00 = R2C1_GT00;
assign R9C1_GT10 = R2C1_GT10;
assign R3C2_GT00 = R2C2_GT00;
assign R3C2_GT10 = R2C2_GT10;
assign R4C2_GT00 = R2C2_GT00;
assign R4C2_GT10 = R2C2_GT10;
assign R5C2_GT00 = R2C2_GT00;
assign R5C2_GT10 = R2C2_GT10;
assign R6C2_GT00 = R2C2_GT00;
assign R6C2_GT10 = R2C2_GT10;
assign R7C2_GT00 = R2C2_GT00;
assign R7C2_GT10 = R2C2_GT10;
assign R8C2_GT00 = R2C2_GT00;
assign R8C2_GT10 = R2C2_GT10;
assign R9C2_GT00 = R2C2_GT00;
assign R9C2_GT10 = R2C2_GT10;
assign R3C3_GT00 = R2C3_GT00;
assign R3C3_GT10 = R2C3_GT10;
assign R4C3_GT00 = R2C3_GT00;
assign R4C3_GT10 = R2C3_GT10;
assign R5C3_GT00 = R2C3_GT00;
assign R5C3_GT10 = R2C3_GT10;
assign R6C3_GT00 = R2C3_GT00;
assign R6C3_GT10 = R2C3_GT10;
assign R7C3_GT00 = R2C3_GT00;
assign R7C3_GT10 = R2C3_GT10;
assign R8C3_GT00 = R2C3_GT00;
assign R8C3_GT10 = R2C3_GT10;
assign R9C3_GT00 = R2C3_GT00;
assign R9C3_GT10 = R2C3_GT10;
assign R3C4_GT00 = R2C4_GT00;
assign R3C4_GT10 = R2C4_GT10;
assign R4C4_GT00 = R2C4_GT00;
assign R4C4_GT10 = R2C4_GT10;
assign R5C4_GT00 = R2C4_GT00;
assign R5C4_GT10 = R2C4_GT10;
assign R6C4_GT00 = R2C4_GT00;
assign R6C4_GT10 = R2C4_GT10;
assign R7C4_GT00 = R2C4_GT00;
assign R7C4_GT10 = R2C4_GT10;
assign R8C4_GT00 = R2C4_GT00;
assign R8C4_GT10 = R2C4_GT10;
assign R9C4_GT00 = R2C4_GT00;
assign R9C4_GT10 = R2C4_GT10;
assign R3C5_GT00 = R2C5_GT00;
assign R3C5_GT10 = R2C5_GT10;
assign R4C5_GT00 = R2C5_GT00;
assign R4C5_GT10 = R2C5_GT10;
assign R5C5_GT00 = R2C5_GT00;
assign R5C5_GT10 = R2C5_GT10;
assign R6C5_GT00 = R2C5_GT00;
assign R6C5_GT10 = R2C5_GT10;
assign R7C5_GT00 = R2C5_GT00;
assign R7C5_GT10 = R2C5_GT10;
assign R8C5_GT00 = R2C5_GT00;
assign R8C5_GT10 = R2C5_GT10;
assign R9C5_GT00 = R2C5_GT00;
assign R9C5_GT10 = R2C5_GT10;
assign R3C6_GT00 = R2C6_GT00;
assign R3C6_GT10 = R2C6_GT10;
assign R4C6_GT00 = R2C6_GT00;
assign R4C6_GT10 = R2C6_GT10;
assign R5C6_GT00 = R2C6_GT00;
assign R5C6_GT10 = R2C6_GT10;
assign R6C6_GT00 = R2C6_GT00;
assign R6C6_GT10 = R2C6_GT10;
assign R7C6_GT00 = R2C6_GT00;
assign R7C6_GT10 = R2C6_GT10;
assign R8C6_GT00 = R2C6_GT00;
assign R8C6_GT10 = R2C6_GT10;
assign R9C6_GT00 = R2C6_GT00;
assign R9C6_GT10 = R2C6_GT10;
assign R3C7_GT00 = R2C7_GT00;
assign R3C7_GT10 = R2C7_GT10;
assign R4C7_GT00 = R2C7_GT00;
assign R4C7_GT10 = R2C7_GT10;
assign R5C7_GT00 = R2C7_GT00;
assign R5C7_GT10 = R2C7_GT10;
assign R6C7_GT00 = R2C7_GT00;
assign R6C7_GT10 = R2C7_GT10;
assign R7C7_GT00 = R2C7_GT00;
assign R7C7_GT10 = R2C7_GT10;
assign R8C7_GT00 = R2C7_GT00;
assign R8C7_GT10 = R2C7_GT10;
assign R9C7_GT00 = R2C7_GT00;
assign R9C7_GT10 = R2C7_GT10;
assign R3C8_GT00 = R2C8_GT00;
assign R3C8_GT10 = R2C8_GT10;
assign R4C8_GT00 = R2C8_GT00;
assign R4C8_GT10 = R2C8_GT10;
assign R5C8_GT00 = R2C8_GT00;
assign R5C8_GT10 = R2C8_GT10;
assign R6C8_GT00 = R2C8_GT00;
assign R6C8_GT10 = R2C8_GT10;
assign R7C8_GT00 = R2C8_GT00;
assign R7C8_GT10 = R2C8_GT10;
assign R8C8_GT00 = R2C8_GT00;
assign R8C8_GT10 = R2C8_GT10;
assign R9C8_GT00 = R2C8_GT00;
assign R9C8_GT10 = R2C8_GT10;
assign R3C9_GT00 = R2C9_GT00;
assign R3C9_GT10 = R2C9_GT10;
assign R4C9_GT00 = R2C9_GT00;
assign R4C9_GT10 = R2C9_GT10;
assign R5C9_GT00 = R2C9_GT00;
assign R5C9_GT10 = R2C9_GT10;
assign R6C9_GT00 = R2C9_GT00;
assign R6C9_GT10 = R2C9_GT10;
assign R7C9_GT00 = R2C9_GT00;
assign R7C9_GT10 = R2C9_GT10;
assign R8C9_GT00 = R2C9_GT00;
assign R8C9_GT10 = R2C9_GT10;
assign R9C9_GT00 = R2C9_GT00;
assign R9C9_GT10 = R2C9_GT10;
assign R3C10_GT00 = R2C10_GT00;
assign R3C10_GT10 = R2C10_GT10;
assign R4C10_GT00 = R2C10_GT00;
assign R4C10_GT10 = R2C10_GT10;
assign R5C10_GT00 = R2C10_GT00;
assign R5C10_GT10 = R2C10_GT10;
assign R6C10_GT00 = R2C10_GT00;
assign R6C10_GT10 = R2C10_GT10;
assign R7C10_GT00 = R2C10_GT00;
assign R7C10_GT10 = R2C10_GT10;
assign R8C10_GT00 = R2C10_GT00;
assign R8C10_GT10 = R2C10_GT10;
assign R9C10_GT00 = R2C10_GT00;
assign R9C10_GT10 = R2C10_GT10;
assign R3C11_GT00 = R2C11_GT00;
assign R3C11_GT10 = R2C11_GT10;
assign R4C11_GT00 = R2C11_GT00;
assign R4C11_GT10 = R2C11_GT10;
assign R5C11_GT00 = R2C11_GT00;
assign R5C11_GT10 = R2C11_GT10;
assign R6C11_GT00 = R2C11_GT00;
assign R6C11_GT10 = R2C11_GT10;
assign R7C11_GT00 = R2C11_GT00;
assign R7C11_GT10 = R2C11_GT10;
assign R8C11_GT00 = R2C11_GT00;
assign R8C11_GT10 = R2C11_GT10;
assign R9C11_GT00 = R2C11_GT00;
assign R9C11_GT10 = R2C11_GT10;
assign R3C12_GT00 = R2C12_GT00;
assign R3C12_GT10 = R2C12_GT10;
assign R4C12_GT00 = R2C12_GT00;
assign R4C12_GT10 = R2C12_GT10;
assign R5C12_GT00 = R2C12_GT00;
assign R5C12_GT10 = R2C12_GT10;
assign R6C12_GT00 = R2C12_GT00;
assign R6C12_GT10 = R2C12_GT10;
assign R7C12_GT00 = R2C12_GT00;
assign R7C12_GT10 = R2C12_GT10;
assign R8C12_GT00 = R2C12_GT00;
assign R8C12_GT10 = R2C12_GT10;
assign R9C12_GT00 = R2C12_GT00;
assign R9C12_GT10 = R2C12_GT10;
assign R3C13_GT00 = R2C13_GT00;
assign R3C13_GT10 = R2C13_GT10;
assign R4C13_GT00 = R2C13_GT00;
assign R4C13_GT10 = R2C13_GT10;
assign R5C13_GT00 = R2C13_GT00;
assign R5C13_GT10 = R2C13_GT10;
assign R6C13_GT00 = R2C13_GT00;
assign R6C13_GT10 = R2C13_GT10;
assign R7C13_GT00 = R2C13_GT00;
assign R7C13_GT10 = R2C13_GT10;
assign R8C13_GT00 = R2C13_GT00;
assign R8C13_GT10 = R2C13_GT10;
assign R9C13_GT00 = R2C13_GT00;
assign R9C13_GT10 = R2C13_GT10;
assign R3C14_GT00 = R2C14_GT00;
assign R3C14_GT10 = R2C14_GT10;
assign R4C14_GT00 = R2C14_GT00;
assign R4C14_GT10 = R2C14_GT10;
assign R5C14_GT00 = R2C14_GT00;
assign R5C14_GT10 = R2C14_GT10;
assign R6C14_GT00 = R2C14_GT00;
assign R6C14_GT10 = R2C14_GT10;
assign R7C14_GT00 = R2C14_GT00;
assign R7C14_GT10 = R2C14_GT10;
assign R8C14_GT00 = R2C14_GT00;
assign R8C14_GT10 = R2C14_GT10;
assign R9C14_GT00 = R2C14_GT00;
assign R9C14_GT10 = R2C14_GT10;
assign R3C15_GT00 = R2C15_GT00;
assign R3C15_GT10 = R2C15_GT10;
assign R4C15_GT00 = R2C15_GT00;
assign R4C15_GT10 = R2C15_GT10;
assign R5C15_GT00 = R2C15_GT00;
assign R5C15_GT10 = R2C15_GT10;
assign R6C15_GT00 = R2C15_GT00;
assign R6C15_GT10 = R2C15_GT10;
assign R7C15_GT00 = R2C15_GT00;
assign R7C15_GT10 = R2C15_GT10;
assign R8C15_GT00 = R2C15_GT00;
assign R8C15_GT10 = R2C15_GT10;
assign R9C15_GT00 = R2C15_GT00;
assign R9C15_GT10 = R2C15_GT10;
assign R3C16_GT00 = R2C16_GT00;
assign R3C16_GT10 = R2C16_GT10;
assign R4C16_GT00 = R2C16_GT00;
assign R4C16_GT10 = R2C16_GT10;
assign R5C16_GT00 = R2C16_GT00;
assign R5C16_GT10 = R2C16_GT10;
assign R6C16_GT00 = R2C16_GT00;
assign R6C16_GT10 = R2C16_GT10;
assign R7C16_GT00 = R2C16_GT00;
assign R7C16_GT10 = R2C16_GT10;
assign R8C16_GT00 = R2C16_GT00;
assign R8C16_GT10 = R2C16_GT10;
assign R9C16_GT00 = R2C16_GT00;
assign R9C16_GT10 = R2C16_GT10;
assign R3C17_GT00 = R2C17_GT00;
assign R3C17_GT10 = R2C17_GT10;
assign R4C17_GT00 = R2C17_GT00;
assign R4C17_GT10 = R2C17_GT10;
assign R5C17_GT00 = R2C17_GT00;
assign R5C17_GT10 = R2C17_GT10;
assign R6C17_GT00 = R2C17_GT00;
assign R6C17_GT10 = R2C17_GT10;
assign R7C17_GT00 = R2C17_GT00;
assign R7C17_GT10 = R2C17_GT10;
assign R8C17_GT00 = R2C17_GT00;
assign R8C17_GT10 = R2C17_GT10;
assign R9C17_GT00 = R2C17_GT00;
assign R9C17_GT10 = R2C17_GT10;
assign R3C18_GT00 = R2C18_GT00;
assign R3C18_GT10 = R2C18_GT10;
assign R4C18_GT00 = R2C18_GT00;
assign R4C18_GT10 = R2C18_GT10;
assign R5C18_GT00 = R2C18_GT00;
assign R5C18_GT10 = R2C18_GT10;
assign R6C18_GT00 = R2C18_GT00;
assign R6C18_GT10 = R2C18_GT10;
assign R7C18_GT00 = R2C18_GT00;
assign R7C18_GT10 = R2C18_GT10;
assign R8C18_GT00 = R2C18_GT00;
assign R8C18_GT10 = R2C18_GT10;
assign R9C18_GT00 = R2C18_GT00;
assign R9C18_GT10 = R2C18_GT10;
assign R3C19_GT00 = R2C19_GT00;
assign R3C19_GT10 = R2C19_GT10;
assign R4C19_GT00 = R2C19_GT00;
assign R4C19_GT10 = R2C19_GT10;
assign R5C19_GT00 = R2C19_GT00;
assign R5C19_GT10 = R2C19_GT10;
assign R6C19_GT00 = R2C19_GT00;
assign R6C19_GT10 = R2C19_GT10;
assign R7C19_GT00 = R2C19_GT00;
assign R7C19_GT10 = R2C19_GT10;
assign R8C19_GT00 = R2C19_GT00;
assign R8C19_GT10 = R2C19_GT10;
assign R9C19_GT00 = R2C19_GT00;
assign R9C19_GT10 = R2C19_GT10;
assign R3C20_GT00 = R2C20_GT00;
assign R3C20_GT10 = R2C20_GT10;
assign R4C20_GT00 = R2C20_GT00;
assign R4C20_GT10 = R2C20_GT10;
assign R5C20_GT00 = R2C20_GT00;
assign R5C20_GT10 = R2C20_GT10;
assign R6C20_GT00 = R2C20_GT00;
assign R6C20_GT10 = R2C20_GT10;
assign R7C20_GT00 = R2C20_GT00;
assign R7C20_GT10 = R2C20_GT10;
assign R8C20_GT00 = R2C20_GT00;
assign R8C20_GT10 = R2C20_GT10;
assign R9C20_GT00 = R2C20_GT00;
assign R9C20_GT10 = R2C20_GT10;
assign R3C21_GT00 = R2C21_GT00;
assign R3C21_GT10 = R2C21_GT10;
assign R4C21_GT00 = R2C21_GT00;
assign R4C21_GT10 = R2C21_GT10;
assign R5C21_GT00 = R2C21_GT00;
assign R5C21_GT10 = R2C21_GT10;
assign R6C21_GT00 = R2C21_GT00;
assign R6C21_GT10 = R2C21_GT10;
assign R7C21_GT00 = R2C21_GT00;
assign R7C21_GT10 = R2C21_GT10;
assign R8C21_GT00 = R2C21_GT00;
assign R8C21_GT10 = R2C21_GT10;
assign R9C21_GT00 = R2C21_GT00;
assign R9C21_GT10 = R2C21_GT10;
assign R3C22_GT00 = R2C22_GT00;
assign R3C22_GT10 = R2C22_GT10;
assign R4C22_GT00 = R2C22_GT00;
assign R4C22_GT10 = R2C22_GT10;
assign R5C22_GT00 = R2C22_GT00;
assign R5C22_GT10 = R2C22_GT10;
assign R6C22_GT00 = R2C22_GT00;
assign R6C22_GT10 = R2C22_GT10;
assign R7C22_GT00 = R2C22_GT00;
assign R7C22_GT10 = R2C22_GT10;
assign R8C22_GT00 = R2C22_GT00;
assign R8C22_GT10 = R2C22_GT10;
assign R9C22_GT00 = R2C22_GT00;
assign R9C22_GT10 = R2C22_GT10;
assign R3C23_GT00 = R2C23_GT00;
assign R3C23_GT10 = R2C23_GT10;
assign R4C23_GT00 = R2C23_GT00;
assign R4C23_GT10 = R2C23_GT10;
assign R5C23_GT00 = R2C23_GT00;
assign R5C23_GT10 = R2C23_GT10;
assign R6C23_GT00 = R2C23_GT00;
assign R6C23_GT10 = R2C23_GT10;
assign R7C23_GT00 = R2C23_GT00;
assign R7C23_GT10 = R2C23_GT10;
assign R8C23_GT00 = R2C23_GT00;
assign R8C23_GT10 = R2C23_GT10;
assign R9C23_GT00 = R2C23_GT00;
assign R9C23_GT10 = R2C23_GT10;
assign R3C24_GT00 = R2C24_GT00;
assign R3C24_GT10 = R2C24_GT10;
assign R4C24_GT00 = R2C24_GT00;
assign R4C24_GT10 = R2C24_GT10;
assign R5C24_GT00 = R2C24_GT00;
assign R5C24_GT10 = R2C24_GT10;
assign R6C24_GT00 = R2C24_GT00;
assign R6C24_GT10 = R2C24_GT10;
assign R7C24_GT00 = R2C24_GT00;
assign R7C24_GT10 = R2C24_GT10;
assign R8C24_GT00 = R2C24_GT00;
assign R8C24_GT10 = R2C24_GT10;
assign R9C24_GT00 = R2C24_GT00;
assign R9C24_GT10 = R2C24_GT10;
assign R3C25_GT00 = R2C25_GT00;
assign R3C25_GT10 = R2C25_GT10;
assign R4C25_GT00 = R2C25_GT00;
assign R4C25_GT10 = R2C25_GT10;
assign R5C25_GT00 = R2C25_GT00;
assign R5C25_GT10 = R2C25_GT10;
assign R6C25_GT00 = R2C25_GT00;
assign R6C25_GT10 = R2C25_GT10;
assign R7C25_GT00 = R2C25_GT00;
assign R7C25_GT10 = R2C25_GT10;
assign R8C25_GT00 = R2C25_GT00;
assign R8C25_GT10 = R2C25_GT10;
assign R9C25_GT00 = R2C25_GT00;
assign R9C25_GT10 = R2C25_GT10;
assign R3C26_GT00 = R2C26_GT00;
assign R3C26_GT10 = R2C26_GT10;
assign R4C26_GT00 = R2C26_GT00;
assign R4C26_GT10 = R2C26_GT10;
assign R5C26_GT00 = R2C26_GT00;
assign R5C26_GT10 = R2C26_GT10;
assign R6C26_GT00 = R2C26_GT00;
assign R6C26_GT10 = R2C26_GT10;
assign R7C26_GT00 = R2C26_GT00;
assign R7C26_GT10 = R2C26_GT10;
assign R8C26_GT00 = R2C26_GT00;
assign R8C26_GT10 = R2C26_GT10;
assign R9C26_GT00 = R2C26_GT00;
assign R9C26_GT10 = R2C26_GT10;
assign R3C27_GT00 = R2C27_GT00;
assign R3C27_GT10 = R2C27_GT10;
assign R4C27_GT00 = R2C27_GT00;
assign R4C27_GT10 = R2C27_GT10;
assign R5C27_GT00 = R2C27_GT00;
assign R5C27_GT10 = R2C27_GT10;
assign R6C27_GT00 = R2C27_GT00;
assign R6C27_GT10 = R2C27_GT10;
assign R7C27_GT00 = R2C27_GT00;
assign R7C27_GT10 = R2C27_GT10;
assign R8C27_GT00 = R2C27_GT00;
assign R8C27_GT10 = R2C27_GT10;
assign R9C27_GT00 = R2C27_GT00;
assign R9C27_GT10 = R2C27_GT10;
assign R3C28_GT00 = R2C28_GT00;
assign R3C28_GT10 = R2C28_GT10;
assign R4C28_GT00 = R2C28_GT00;
assign R4C28_GT10 = R2C28_GT10;
assign R5C28_GT00 = R2C28_GT00;
assign R5C28_GT10 = R2C28_GT10;
assign R6C28_GT00 = R2C28_GT00;
assign R6C28_GT10 = R2C28_GT10;
assign R7C28_GT00 = R2C28_GT00;
assign R7C28_GT10 = R2C28_GT10;
assign R8C28_GT00 = R2C28_GT00;
assign R8C28_GT10 = R2C28_GT10;
assign R9C28_GT00 = R2C28_GT00;
assign R9C28_GT10 = R2C28_GT10;
assign R11C1_GT00 = R20C1_GT00;
assign R11C1_GT10 = R20C1_GT10;
assign R12C1_GT00 = R20C1_GT00;
assign R12C1_GT10 = R20C1_GT10;
assign R13C1_GT00 = R20C1_GT00;
assign R13C1_GT10 = R20C1_GT10;
assign R14C1_GT00 = R20C1_GT00;
assign R14C1_GT10 = R20C1_GT10;
assign R15C1_GT00 = R20C1_GT00;
assign R15C1_GT10 = R20C1_GT10;
assign R16C1_GT00 = R20C1_GT00;
assign R16C1_GT10 = R20C1_GT10;
assign R17C1_GT00 = R20C1_GT00;
assign R17C1_GT10 = R20C1_GT10;
assign R18C1_GT00 = R20C1_GT00;
assign R18C1_GT10 = R20C1_GT10;
assign R21C1_GT00 = R20C1_GT00;
assign R21C1_GT10 = R20C1_GT10;
assign R22C1_GT00 = R20C1_GT00;
assign R22C1_GT10 = R20C1_GT10;
assign R23C1_GT00 = R20C1_GT00;
assign R23C1_GT10 = R20C1_GT10;
assign R24C1_GT00 = R20C1_GT00;
assign R24C1_GT10 = R20C1_GT10;
assign R25C1_GT00 = R20C1_GT00;
assign R25C1_GT10 = R20C1_GT10;
assign R26C1_GT00 = R20C1_GT00;
assign R26C1_GT10 = R20C1_GT10;
assign R27C1_GT00 = R20C1_GT00;
assign R27C1_GT10 = R20C1_GT10;
assign R11C2_GT00 = R20C2_GT00;
assign R11C2_GT10 = R20C2_GT10;
assign R12C2_GT00 = R20C2_GT00;
assign R12C2_GT10 = R20C2_GT10;
assign R13C2_GT00 = R20C2_GT00;
assign R13C2_GT10 = R20C2_GT10;
assign R14C2_GT00 = R20C2_GT00;
assign R14C2_GT10 = R20C2_GT10;
assign R15C2_GT00 = R20C2_GT00;
assign R15C2_GT10 = R20C2_GT10;
assign R16C2_GT00 = R20C2_GT00;
assign R16C2_GT10 = R20C2_GT10;
assign R17C2_GT00 = R20C2_GT00;
assign R17C2_GT10 = R20C2_GT10;
assign R18C2_GT00 = R20C2_GT00;
assign R18C2_GT10 = R20C2_GT10;
assign R21C2_GT00 = R20C2_GT00;
assign R21C2_GT10 = R20C2_GT10;
assign R22C2_GT00 = R20C2_GT00;
assign R22C2_GT10 = R20C2_GT10;
assign R23C2_GT00 = R20C2_GT00;
assign R23C2_GT10 = R20C2_GT10;
assign R24C2_GT00 = R20C2_GT00;
assign R24C2_GT10 = R20C2_GT10;
assign R25C2_GT00 = R20C2_GT00;
assign R25C2_GT10 = R20C2_GT10;
assign R26C2_GT00 = R20C2_GT00;
assign R26C2_GT10 = R20C2_GT10;
assign R27C2_GT00 = R20C2_GT00;
assign R27C2_GT10 = R20C2_GT10;
assign R11C3_GT00 = R20C3_GT00;
assign R11C3_GT10 = R20C3_GT10;
assign R12C3_GT00 = R20C3_GT00;
assign R12C3_GT10 = R20C3_GT10;
assign R13C3_GT00 = R20C3_GT00;
assign R13C3_GT10 = R20C3_GT10;
assign R14C3_GT00 = R20C3_GT00;
assign R14C3_GT10 = R20C3_GT10;
assign R15C3_GT00 = R20C3_GT00;
assign R15C3_GT10 = R20C3_GT10;
assign R16C3_GT00 = R20C3_GT00;
assign R16C3_GT10 = R20C3_GT10;
assign R17C3_GT00 = R20C3_GT00;
assign R17C3_GT10 = R20C3_GT10;
assign R18C3_GT00 = R20C3_GT00;
assign R18C3_GT10 = R20C3_GT10;
assign R21C3_GT00 = R20C3_GT00;
assign R21C3_GT10 = R20C3_GT10;
assign R22C3_GT00 = R20C3_GT00;
assign R22C3_GT10 = R20C3_GT10;
assign R23C3_GT00 = R20C3_GT00;
assign R23C3_GT10 = R20C3_GT10;
assign R24C3_GT00 = R20C3_GT00;
assign R24C3_GT10 = R20C3_GT10;
assign R25C3_GT00 = R20C3_GT00;
assign R25C3_GT10 = R20C3_GT10;
assign R26C3_GT00 = R20C3_GT00;
assign R26C3_GT10 = R20C3_GT10;
assign R27C3_GT00 = R20C3_GT00;
assign R27C3_GT10 = R20C3_GT10;
assign R11C4_GT00 = R20C4_GT00;
assign R11C4_GT10 = R20C4_GT10;
assign R12C4_GT00 = R20C4_GT00;
assign R12C4_GT10 = R20C4_GT10;
assign R13C4_GT00 = R20C4_GT00;
assign R13C4_GT10 = R20C4_GT10;
assign R14C4_GT00 = R20C4_GT00;
assign R14C4_GT10 = R20C4_GT10;
assign R15C4_GT00 = R20C4_GT00;
assign R15C4_GT10 = R20C4_GT10;
assign R16C4_GT00 = R20C4_GT00;
assign R16C4_GT10 = R20C4_GT10;
assign R17C4_GT00 = R20C4_GT00;
assign R17C4_GT10 = R20C4_GT10;
assign R18C4_GT00 = R20C4_GT00;
assign R18C4_GT10 = R20C4_GT10;
assign R21C4_GT00 = R20C4_GT00;
assign R21C4_GT10 = R20C4_GT10;
assign R22C4_GT00 = R20C4_GT00;
assign R22C4_GT10 = R20C4_GT10;
assign R23C4_GT00 = R20C4_GT00;
assign R23C4_GT10 = R20C4_GT10;
assign R24C4_GT00 = R20C4_GT00;
assign R24C4_GT10 = R20C4_GT10;
assign R25C4_GT00 = R20C4_GT00;
assign R25C4_GT10 = R20C4_GT10;
assign R26C4_GT00 = R20C4_GT00;
assign R26C4_GT10 = R20C4_GT10;
assign R27C4_GT00 = R20C4_GT00;
assign R27C4_GT10 = R20C4_GT10;
assign R11C5_GT00 = R20C5_GT00;
assign R11C5_GT10 = R20C5_GT10;
assign R12C5_GT00 = R20C5_GT00;
assign R12C5_GT10 = R20C5_GT10;
assign R13C5_GT00 = R20C5_GT00;
assign R13C5_GT10 = R20C5_GT10;
assign R14C5_GT00 = R20C5_GT00;
assign R14C5_GT10 = R20C5_GT10;
assign R15C5_GT00 = R20C5_GT00;
assign R15C5_GT10 = R20C5_GT10;
assign R16C5_GT00 = R20C5_GT00;
assign R16C5_GT10 = R20C5_GT10;
assign R17C5_GT00 = R20C5_GT00;
assign R17C5_GT10 = R20C5_GT10;
assign R18C5_GT00 = R20C5_GT00;
assign R18C5_GT10 = R20C5_GT10;
assign R21C5_GT00 = R20C5_GT00;
assign R21C5_GT10 = R20C5_GT10;
assign R22C5_GT00 = R20C5_GT00;
assign R22C5_GT10 = R20C5_GT10;
assign R23C5_GT00 = R20C5_GT00;
assign R23C5_GT10 = R20C5_GT10;
assign R24C5_GT00 = R20C5_GT00;
assign R24C5_GT10 = R20C5_GT10;
assign R25C5_GT00 = R20C5_GT00;
assign R25C5_GT10 = R20C5_GT10;
assign R26C5_GT00 = R20C5_GT00;
assign R26C5_GT10 = R20C5_GT10;
assign R27C5_GT00 = R20C5_GT00;
assign R27C5_GT10 = R20C5_GT10;
assign R11C6_GT00 = R20C6_GT00;
assign R11C6_GT10 = R20C6_GT10;
assign R12C6_GT00 = R20C6_GT00;
assign R12C6_GT10 = R20C6_GT10;
assign R13C6_GT00 = R20C6_GT00;
assign R13C6_GT10 = R20C6_GT10;
assign R14C6_GT00 = R20C6_GT00;
assign R14C6_GT10 = R20C6_GT10;
assign R15C6_GT00 = R20C6_GT00;
assign R15C6_GT10 = R20C6_GT10;
assign R16C6_GT00 = R20C6_GT00;
assign R16C6_GT10 = R20C6_GT10;
assign R17C6_GT00 = R20C6_GT00;
assign R17C6_GT10 = R20C6_GT10;
assign R18C6_GT00 = R20C6_GT00;
assign R18C6_GT10 = R20C6_GT10;
assign R21C6_GT00 = R20C6_GT00;
assign R21C6_GT10 = R20C6_GT10;
assign R22C6_GT00 = R20C6_GT00;
assign R22C6_GT10 = R20C6_GT10;
assign R23C6_GT00 = R20C6_GT00;
assign R23C6_GT10 = R20C6_GT10;
assign R24C6_GT00 = R20C6_GT00;
assign R24C6_GT10 = R20C6_GT10;
assign R25C6_GT00 = R20C6_GT00;
assign R25C6_GT10 = R20C6_GT10;
assign R26C6_GT00 = R20C6_GT00;
assign R26C6_GT10 = R20C6_GT10;
assign R27C6_GT00 = R20C6_GT00;
assign R27C6_GT10 = R20C6_GT10;
assign R11C7_GT00 = R20C7_GT00;
assign R11C7_GT10 = R20C7_GT10;
assign R12C7_GT00 = R20C7_GT00;
assign R12C7_GT10 = R20C7_GT10;
assign R13C7_GT00 = R20C7_GT00;
assign R13C7_GT10 = R20C7_GT10;
assign R14C7_GT00 = R20C7_GT00;
assign R14C7_GT10 = R20C7_GT10;
assign R15C7_GT00 = R20C7_GT00;
assign R15C7_GT10 = R20C7_GT10;
assign R16C7_GT00 = R20C7_GT00;
assign R16C7_GT10 = R20C7_GT10;
assign R17C7_GT00 = R20C7_GT00;
assign R17C7_GT10 = R20C7_GT10;
assign R18C7_GT00 = R20C7_GT00;
assign R18C7_GT10 = R20C7_GT10;
assign R21C7_GT00 = R20C7_GT00;
assign R21C7_GT10 = R20C7_GT10;
assign R22C7_GT00 = R20C7_GT00;
assign R22C7_GT10 = R20C7_GT10;
assign R23C7_GT00 = R20C7_GT00;
assign R23C7_GT10 = R20C7_GT10;
assign R24C7_GT00 = R20C7_GT00;
assign R24C7_GT10 = R20C7_GT10;
assign R25C7_GT00 = R20C7_GT00;
assign R25C7_GT10 = R20C7_GT10;
assign R26C7_GT00 = R20C7_GT00;
assign R26C7_GT10 = R20C7_GT10;
assign R27C7_GT00 = R20C7_GT00;
assign R27C7_GT10 = R20C7_GT10;
assign R11C8_GT00 = R20C8_GT00;
assign R11C8_GT10 = R20C8_GT10;
assign R12C8_GT00 = R20C8_GT00;
assign R12C8_GT10 = R20C8_GT10;
assign R13C8_GT00 = R20C8_GT00;
assign R13C8_GT10 = R20C8_GT10;
assign R14C8_GT00 = R20C8_GT00;
assign R14C8_GT10 = R20C8_GT10;
assign R15C8_GT00 = R20C8_GT00;
assign R15C8_GT10 = R20C8_GT10;
assign R16C8_GT00 = R20C8_GT00;
assign R16C8_GT10 = R20C8_GT10;
assign R17C8_GT00 = R20C8_GT00;
assign R17C8_GT10 = R20C8_GT10;
assign R18C8_GT00 = R20C8_GT00;
assign R18C8_GT10 = R20C8_GT10;
assign R21C8_GT00 = R20C8_GT00;
assign R21C8_GT10 = R20C8_GT10;
assign R22C8_GT00 = R20C8_GT00;
assign R22C8_GT10 = R20C8_GT10;
assign R23C8_GT00 = R20C8_GT00;
assign R23C8_GT10 = R20C8_GT10;
assign R24C8_GT00 = R20C8_GT00;
assign R24C8_GT10 = R20C8_GT10;
assign R25C8_GT00 = R20C8_GT00;
assign R25C8_GT10 = R20C8_GT10;
assign R26C8_GT00 = R20C8_GT00;
assign R26C8_GT10 = R20C8_GT10;
assign R27C8_GT00 = R20C8_GT00;
assign R27C8_GT10 = R20C8_GT10;
assign R11C9_GT00 = R20C9_GT00;
assign R11C9_GT10 = R20C9_GT10;
assign R12C9_GT00 = R20C9_GT00;
assign R12C9_GT10 = R20C9_GT10;
assign R13C9_GT00 = R20C9_GT00;
assign R13C9_GT10 = R20C9_GT10;
assign R14C9_GT00 = R20C9_GT00;
assign R14C9_GT10 = R20C9_GT10;
assign R15C9_GT00 = R20C9_GT00;
assign R15C9_GT10 = R20C9_GT10;
assign R16C9_GT00 = R20C9_GT00;
assign R16C9_GT10 = R20C9_GT10;
assign R17C9_GT00 = R20C9_GT00;
assign R17C9_GT10 = R20C9_GT10;
assign R18C9_GT00 = R20C9_GT00;
assign R18C9_GT10 = R20C9_GT10;
assign R21C9_GT00 = R20C9_GT00;
assign R21C9_GT10 = R20C9_GT10;
assign R22C9_GT00 = R20C9_GT00;
assign R22C9_GT10 = R20C9_GT10;
assign R23C9_GT00 = R20C9_GT00;
assign R23C9_GT10 = R20C9_GT10;
assign R24C9_GT00 = R20C9_GT00;
assign R24C9_GT10 = R20C9_GT10;
assign R25C9_GT00 = R20C9_GT00;
assign R25C9_GT10 = R20C9_GT10;
assign R26C9_GT00 = R20C9_GT00;
assign R26C9_GT10 = R20C9_GT10;
assign R27C9_GT00 = R20C9_GT00;
assign R27C9_GT10 = R20C9_GT10;
assign R11C10_GT00 = R20C10_GT00;
assign R11C10_GT10 = R20C10_GT10;
assign R12C10_GT00 = R20C10_GT00;
assign R12C10_GT10 = R20C10_GT10;
assign R13C10_GT00 = R20C10_GT00;
assign R13C10_GT10 = R20C10_GT10;
assign R14C10_GT00 = R20C10_GT00;
assign R14C10_GT10 = R20C10_GT10;
assign R15C10_GT00 = R20C10_GT00;
assign R15C10_GT10 = R20C10_GT10;
assign R16C10_GT00 = R20C10_GT00;
assign R16C10_GT10 = R20C10_GT10;
assign R17C10_GT00 = R20C10_GT00;
assign R17C10_GT10 = R20C10_GT10;
assign R18C10_GT00 = R20C10_GT00;
assign R18C10_GT10 = R20C10_GT10;
assign R21C10_GT00 = R20C10_GT00;
assign R21C10_GT10 = R20C10_GT10;
assign R22C10_GT00 = R20C10_GT00;
assign R22C10_GT10 = R20C10_GT10;
assign R23C10_GT00 = R20C10_GT00;
assign R23C10_GT10 = R20C10_GT10;
assign R24C10_GT00 = R20C10_GT00;
assign R24C10_GT10 = R20C10_GT10;
assign R25C10_GT00 = R20C10_GT00;
assign R25C10_GT10 = R20C10_GT10;
assign R26C10_GT00 = R20C10_GT00;
assign R26C10_GT10 = R20C10_GT10;
assign R27C10_GT00 = R20C10_GT00;
assign R27C10_GT10 = R20C10_GT10;
assign R11C11_GT00 = R20C11_GT00;
assign R11C11_GT10 = R20C11_GT10;
assign R12C11_GT00 = R20C11_GT00;
assign R12C11_GT10 = R20C11_GT10;
assign R13C11_GT00 = R20C11_GT00;
assign R13C11_GT10 = R20C11_GT10;
assign R14C11_GT00 = R20C11_GT00;
assign R14C11_GT10 = R20C11_GT10;
assign R15C11_GT00 = R20C11_GT00;
assign R15C11_GT10 = R20C11_GT10;
assign R16C11_GT00 = R20C11_GT00;
assign R16C11_GT10 = R20C11_GT10;
assign R17C11_GT00 = R20C11_GT00;
assign R17C11_GT10 = R20C11_GT10;
assign R18C11_GT00 = R20C11_GT00;
assign R18C11_GT10 = R20C11_GT10;
assign R21C11_GT00 = R20C11_GT00;
assign R21C11_GT10 = R20C11_GT10;
assign R22C11_GT00 = R20C11_GT00;
assign R22C11_GT10 = R20C11_GT10;
assign R23C11_GT00 = R20C11_GT00;
assign R23C11_GT10 = R20C11_GT10;
assign R24C11_GT00 = R20C11_GT00;
assign R24C11_GT10 = R20C11_GT10;
assign R25C11_GT00 = R20C11_GT00;
assign R25C11_GT10 = R20C11_GT10;
assign R26C11_GT00 = R20C11_GT00;
assign R26C11_GT10 = R20C11_GT10;
assign R27C11_GT00 = R20C11_GT00;
assign R27C11_GT10 = R20C11_GT10;
assign R11C12_GT00 = R20C12_GT00;
assign R11C12_GT10 = R20C12_GT10;
assign R12C12_GT00 = R20C12_GT00;
assign R12C12_GT10 = R20C12_GT10;
assign R13C12_GT00 = R20C12_GT00;
assign R13C12_GT10 = R20C12_GT10;
assign R14C12_GT00 = R20C12_GT00;
assign R14C12_GT10 = R20C12_GT10;
assign R15C12_GT00 = R20C12_GT00;
assign R15C12_GT10 = R20C12_GT10;
assign R16C12_GT00 = R20C12_GT00;
assign R16C12_GT10 = R20C12_GT10;
assign R17C12_GT00 = R20C12_GT00;
assign R17C12_GT10 = R20C12_GT10;
assign R18C12_GT00 = R20C12_GT00;
assign R18C12_GT10 = R20C12_GT10;
assign R21C12_GT00 = R20C12_GT00;
assign R21C12_GT10 = R20C12_GT10;
assign R22C12_GT00 = R20C12_GT00;
assign R22C12_GT10 = R20C12_GT10;
assign R23C12_GT00 = R20C12_GT00;
assign R23C12_GT10 = R20C12_GT10;
assign R24C12_GT00 = R20C12_GT00;
assign R24C12_GT10 = R20C12_GT10;
assign R25C12_GT00 = R20C12_GT00;
assign R25C12_GT10 = R20C12_GT10;
assign R26C12_GT00 = R20C12_GT00;
assign R26C12_GT10 = R20C12_GT10;
assign R27C12_GT00 = R20C12_GT00;
assign R27C12_GT10 = R20C12_GT10;
assign R11C13_GT00 = R20C13_GT00;
assign R11C13_GT10 = R20C13_GT10;
assign R12C13_GT00 = R20C13_GT00;
assign R12C13_GT10 = R20C13_GT10;
assign R13C13_GT00 = R20C13_GT00;
assign R13C13_GT10 = R20C13_GT10;
assign R14C13_GT00 = R20C13_GT00;
assign R14C13_GT10 = R20C13_GT10;
assign R15C13_GT00 = R20C13_GT00;
assign R15C13_GT10 = R20C13_GT10;
assign R16C13_GT00 = R20C13_GT00;
assign R16C13_GT10 = R20C13_GT10;
assign R17C13_GT00 = R20C13_GT00;
assign R17C13_GT10 = R20C13_GT10;
assign R18C13_GT00 = R20C13_GT00;
assign R18C13_GT10 = R20C13_GT10;
assign R21C13_GT00 = R20C13_GT00;
assign R21C13_GT10 = R20C13_GT10;
assign R22C13_GT00 = R20C13_GT00;
assign R22C13_GT10 = R20C13_GT10;
assign R23C13_GT00 = R20C13_GT00;
assign R23C13_GT10 = R20C13_GT10;
assign R24C13_GT00 = R20C13_GT00;
assign R24C13_GT10 = R20C13_GT10;
assign R25C13_GT00 = R20C13_GT00;
assign R25C13_GT10 = R20C13_GT10;
assign R26C13_GT00 = R20C13_GT00;
assign R26C13_GT10 = R20C13_GT10;
assign R27C13_GT00 = R20C13_GT00;
assign R27C13_GT10 = R20C13_GT10;
assign R11C14_GT00 = R20C14_GT00;
assign R11C14_GT10 = R20C14_GT10;
assign R12C14_GT00 = R20C14_GT00;
assign R12C14_GT10 = R20C14_GT10;
assign R13C14_GT00 = R20C14_GT00;
assign R13C14_GT10 = R20C14_GT10;
assign R14C14_GT00 = R20C14_GT00;
assign R14C14_GT10 = R20C14_GT10;
assign R15C14_GT00 = R20C14_GT00;
assign R15C14_GT10 = R20C14_GT10;
assign R16C14_GT00 = R20C14_GT00;
assign R16C14_GT10 = R20C14_GT10;
assign R17C14_GT00 = R20C14_GT00;
assign R17C14_GT10 = R20C14_GT10;
assign R18C14_GT00 = R20C14_GT00;
assign R18C14_GT10 = R20C14_GT10;
assign R21C14_GT00 = R20C14_GT00;
assign R21C14_GT10 = R20C14_GT10;
assign R22C14_GT00 = R20C14_GT00;
assign R22C14_GT10 = R20C14_GT10;
assign R23C14_GT00 = R20C14_GT00;
assign R23C14_GT10 = R20C14_GT10;
assign R24C14_GT00 = R20C14_GT00;
assign R24C14_GT10 = R20C14_GT10;
assign R25C14_GT00 = R20C14_GT00;
assign R25C14_GT10 = R20C14_GT10;
assign R26C14_GT00 = R20C14_GT00;
assign R26C14_GT10 = R20C14_GT10;
assign R27C14_GT00 = R20C14_GT00;
assign R27C14_GT10 = R20C14_GT10;
assign R11C15_GT00 = R20C15_GT00;
assign R11C15_GT10 = R20C15_GT10;
assign R12C15_GT00 = R20C15_GT00;
assign R12C15_GT10 = R20C15_GT10;
assign R13C15_GT00 = R20C15_GT00;
assign R13C15_GT10 = R20C15_GT10;
assign R14C15_GT00 = R20C15_GT00;
assign R14C15_GT10 = R20C15_GT10;
assign R15C15_GT00 = R20C15_GT00;
assign R15C15_GT10 = R20C15_GT10;
assign R16C15_GT00 = R20C15_GT00;
assign R16C15_GT10 = R20C15_GT10;
assign R17C15_GT00 = R20C15_GT00;
assign R17C15_GT10 = R20C15_GT10;
assign R18C15_GT00 = R20C15_GT00;
assign R18C15_GT10 = R20C15_GT10;
assign R21C15_GT00 = R20C15_GT00;
assign R21C15_GT10 = R20C15_GT10;
assign R22C15_GT00 = R20C15_GT00;
assign R22C15_GT10 = R20C15_GT10;
assign R23C15_GT00 = R20C15_GT00;
assign R23C15_GT10 = R20C15_GT10;
assign R24C15_GT00 = R20C15_GT00;
assign R24C15_GT10 = R20C15_GT10;
assign R25C15_GT00 = R20C15_GT00;
assign R25C15_GT10 = R20C15_GT10;
assign R26C15_GT00 = R20C15_GT00;
assign R26C15_GT10 = R20C15_GT10;
assign R27C15_GT00 = R20C15_GT00;
assign R27C15_GT10 = R20C15_GT10;
assign R11C16_GT00 = R20C16_GT00;
assign R11C16_GT10 = R20C16_GT10;
assign R12C16_GT00 = R20C16_GT00;
assign R12C16_GT10 = R20C16_GT10;
assign R13C16_GT00 = R20C16_GT00;
assign R13C16_GT10 = R20C16_GT10;
assign R14C16_GT00 = R20C16_GT00;
assign R14C16_GT10 = R20C16_GT10;
assign R15C16_GT00 = R20C16_GT00;
assign R15C16_GT10 = R20C16_GT10;
assign R16C16_GT00 = R20C16_GT00;
assign R16C16_GT10 = R20C16_GT10;
assign R17C16_GT00 = R20C16_GT00;
assign R17C16_GT10 = R20C16_GT10;
assign R18C16_GT00 = R20C16_GT00;
assign R18C16_GT10 = R20C16_GT10;
assign R21C16_GT00 = R20C16_GT00;
assign R21C16_GT10 = R20C16_GT10;
assign R22C16_GT00 = R20C16_GT00;
assign R22C16_GT10 = R20C16_GT10;
assign R23C16_GT00 = R20C16_GT00;
assign R23C16_GT10 = R20C16_GT10;
assign R24C16_GT00 = R20C16_GT00;
assign R24C16_GT10 = R20C16_GT10;
assign R25C16_GT00 = R20C16_GT00;
assign R25C16_GT10 = R20C16_GT10;
assign R26C16_GT00 = R20C16_GT00;
assign R26C16_GT10 = R20C16_GT10;
assign R27C16_GT00 = R20C16_GT00;
assign R27C16_GT10 = R20C16_GT10;
assign R11C17_GT00 = R20C17_GT00;
assign R11C17_GT10 = R20C17_GT10;
assign R12C17_GT00 = R20C17_GT00;
assign R12C17_GT10 = R20C17_GT10;
assign R13C17_GT00 = R20C17_GT00;
assign R13C17_GT10 = R20C17_GT10;
assign R14C17_GT00 = R20C17_GT00;
assign R14C17_GT10 = R20C17_GT10;
assign R15C17_GT00 = R20C17_GT00;
assign R15C17_GT10 = R20C17_GT10;
assign R16C17_GT00 = R20C17_GT00;
assign R16C17_GT10 = R20C17_GT10;
assign R17C17_GT00 = R20C17_GT00;
assign R17C17_GT10 = R20C17_GT10;
assign R18C17_GT00 = R20C17_GT00;
assign R18C17_GT10 = R20C17_GT10;
assign R21C17_GT00 = R20C17_GT00;
assign R21C17_GT10 = R20C17_GT10;
assign R22C17_GT00 = R20C17_GT00;
assign R22C17_GT10 = R20C17_GT10;
assign R23C17_GT00 = R20C17_GT00;
assign R23C17_GT10 = R20C17_GT10;
assign R24C17_GT00 = R20C17_GT00;
assign R24C17_GT10 = R20C17_GT10;
assign R25C17_GT00 = R20C17_GT00;
assign R25C17_GT10 = R20C17_GT10;
assign R26C17_GT00 = R20C17_GT00;
assign R26C17_GT10 = R20C17_GT10;
assign R27C17_GT00 = R20C17_GT00;
assign R27C17_GT10 = R20C17_GT10;
assign R11C18_GT00 = R20C18_GT00;
assign R11C18_GT10 = R20C18_GT10;
assign R12C18_GT00 = R20C18_GT00;
assign R12C18_GT10 = R20C18_GT10;
assign R13C18_GT00 = R20C18_GT00;
assign R13C18_GT10 = R20C18_GT10;
assign R14C18_GT00 = R20C18_GT00;
assign R14C18_GT10 = R20C18_GT10;
assign R15C18_GT00 = R20C18_GT00;
assign R15C18_GT10 = R20C18_GT10;
assign R16C18_GT00 = R20C18_GT00;
assign R16C18_GT10 = R20C18_GT10;
assign R17C18_GT00 = R20C18_GT00;
assign R17C18_GT10 = R20C18_GT10;
assign R18C18_GT00 = R20C18_GT00;
assign R18C18_GT10 = R20C18_GT10;
assign R21C18_GT00 = R20C18_GT00;
assign R21C18_GT10 = R20C18_GT10;
assign R22C18_GT00 = R20C18_GT00;
assign R22C18_GT10 = R20C18_GT10;
assign R23C18_GT00 = R20C18_GT00;
assign R23C18_GT10 = R20C18_GT10;
assign R24C18_GT00 = R20C18_GT00;
assign R24C18_GT10 = R20C18_GT10;
assign R25C18_GT00 = R20C18_GT00;
assign R25C18_GT10 = R20C18_GT10;
assign R26C18_GT00 = R20C18_GT00;
assign R26C18_GT10 = R20C18_GT10;
assign R27C18_GT00 = R20C18_GT00;
assign R27C18_GT10 = R20C18_GT10;
assign R11C19_GT00 = R20C19_GT00;
assign R11C19_GT10 = R20C19_GT10;
assign R12C19_GT00 = R20C19_GT00;
assign R12C19_GT10 = R20C19_GT10;
assign R13C19_GT00 = R20C19_GT00;
assign R13C19_GT10 = R20C19_GT10;
assign R14C19_GT00 = R20C19_GT00;
assign R14C19_GT10 = R20C19_GT10;
assign R15C19_GT00 = R20C19_GT00;
assign R15C19_GT10 = R20C19_GT10;
assign R16C19_GT00 = R20C19_GT00;
assign R16C19_GT10 = R20C19_GT10;
assign R17C19_GT00 = R20C19_GT00;
assign R17C19_GT10 = R20C19_GT10;
assign R18C19_GT00 = R20C19_GT00;
assign R18C19_GT10 = R20C19_GT10;
assign R21C19_GT00 = R20C19_GT00;
assign R21C19_GT10 = R20C19_GT10;
assign R22C19_GT00 = R20C19_GT00;
assign R22C19_GT10 = R20C19_GT10;
assign R23C19_GT00 = R20C19_GT00;
assign R23C19_GT10 = R20C19_GT10;
assign R24C19_GT00 = R20C19_GT00;
assign R24C19_GT10 = R20C19_GT10;
assign R25C19_GT00 = R20C19_GT00;
assign R25C19_GT10 = R20C19_GT10;
assign R26C19_GT00 = R20C19_GT00;
assign R26C19_GT10 = R20C19_GT10;
assign R27C19_GT00 = R20C19_GT00;
assign R27C19_GT10 = R20C19_GT10;
assign R11C20_GT00 = R20C20_GT00;
assign R11C20_GT10 = R20C20_GT10;
assign R12C20_GT00 = R20C20_GT00;
assign R12C20_GT10 = R20C20_GT10;
assign R13C20_GT00 = R20C20_GT00;
assign R13C20_GT10 = R20C20_GT10;
assign R14C20_GT00 = R20C20_GT00;
assign R14C20_GT10 = R20C20_GT10;
assign R15C20_GT00 = R20C20_GT00;
assign R15C20_GT10 = R20C20_GT10;
assign R16C20_GT00 = R20C20_GT00;
assign R16C20_GT10 = R20C20_GT10;
assign R17C20_GT00 = R20C20_GT00;
assign R17C20_GT10 = R20C20_GT10;
assign R18C20_GT00 = R20C20_GT00;
assign R18C20_GT10 = R20C20_GT10;
assign R21C20_GT00 = R20C20_GT00;
assign R21C20_GT10 = R20C20_GT10;
assign R22C20_GT00 = R20C20_GT00;
assign R22C20_GT10 = R20C20_GT10;
assign R23C20_GT00 = R20C20_GT00;
assign R23C20_GT10 = R20C20_GT10;
assign R24C20_GT00 = R20C20_GT00;
assign R24C20_GT10 = R20C20_GT10;
assign R25C20_GT00 = R20C20_GT00;
assign R25C20_GT10 = R20C20_GT10;
assign R26C20_GT00 = R20C20_GT00;
assign R26C20_GT10 = R20C20_GT10;
assign R27C20_GT00 = R20C20_GT00;
assign R27C20_GT10 = R20C20_GT10;
assign R11C21_GT00 = R20C21_GT00;
assign R11C21_GT10 = R20C21_GT10;
assign R12C21_GT00 = R20C21_GT00;
assign R12C21_GT10 = R20C21_GT10;
assign R13C21_GT00 = R20C21_GT00;
assign R13C21_GT10 = R20C21_GT10;
assign R14C21_GT00 = R20C21_GT00;
assign R14C21_GT10 = R20C21_GT10;
assign R15C21_GT00 = R20C21_GT00;
assign R15C21_GT10 = R20C21_GT10;
assign R16C21_GT00 = R20C21_GT00;
assign R16C21_GT10 = R20C21_GT10;
assign R17C21_GT00 = R20C21_GT00;
assign R17C21_GT10 = R20C21_GT10;
assign R18C21_GT00 = R20C21_GT00;
assign R18C21_GT10 = R20C21_GT10;
assign R21C21_GT00 = R20C21_GT00;
assign R21C21_GT10 = R20C21_GT10;
assign R22C21_GT00 = R20C21_GT00;
assign R22C21_GT10 = R20C21_GT10;
assign R23C21_GT00 = R20C21_GT00;
assign R23C21_GT10 = R20C21_GT10;
assign R24C21_GT00 = R20C21_GT00;
assign R24C21_GT10 = R20C21_GT10;
assign R25C21_GT00 = R20C21_GT00;
assign R25C21_GT10 = R20C21_GT10;
assign R26C21_GT00 = R20C21_GT00;
assign R26C21_GT10 = R20C21_GT10;
assign R27C21_GT00 = R20C21_GT00;
assign R27C21_GT10 = R20C21_GT10;
assign R11C22_GT00 = R20C22_GT00;
assign R11C22_GT10 = R20C22_GT10;
assign R12C22_GT00 = R20C22_GT00;
assign R12C22_GT10 = R20C22_GT10;
assign R13C22_GT00 = R20C22_GT00;
assign R13C22_GT10 = R20C22_GT10;
assign R14C22_GT00 = R20C22_GT00;
assign R14C22_GT10 = R20C22_GT10;
assign R15C22_GT00 = R20C22_GT00;
assign R15C22_GT10 = R20C22_GT10;
assign R16C22_GT00 = R20C22_GT00;
assign R16C22_GT10 = R20C22_GT10;
assign R17C22_GT00 = R20C22_GT00;
assign R17C22_GT10 = R20C22_GT10;
assign R18C22_GT00 = R20C22_GT00;
assign R18C22_GT10 = R20C22_GT10;
assign R21C22_GT00 = R20C22_GT00;
assign R21C22_GT10 = R20C22_GT10;
assign R22C22_GT00 = R20C22_GT00;
assign R22C22_GT10 = R20C22_GT10;
assign R23C22_GT00 = R20C22_GT00;
assign R23C22_GT10 = R20C22_GT10;
assign R24C22_GT00 = R20C22_GT00;
assign R24C22_GT10 = R20C22_GT10;
assign R25C22_GT00 = R20C22_GT00;
assign R25C22_GT10 = R20C22_GT10;
assign R26C22_GT00 = R20C22_GT00;
assign R26C22_GT10 = R20C22_GT10;
assign R27C22_GT00 = R20C22_GT00;
assign R27C22_GT10 = R20C22_GT10;
assign R11C23_GT00 = R20C23_GT00;
assign R11C23_GT10 = R20C23_GT10;
assign R12C23_GT00 = R20C23_GT00;
assign R12C23_GT10 = R20C23_GT10;
assign R13C23_GT00 = R20C23_GT00;
assign R13C23_GT10 = R20C23_GT10;
assign R14C23_GT00 = R20C23_GT00;
assign R14C23_GT10 = R20C23_GT10;
assign R15C23_GT00 = R20C23_GT00;
assign R15C23_GT10 = R20C23_GT10;
assign R16C23_GT00 = R20C23_GT00;
assign R16C23_GT10 = R20C23_GT10;
assign R17C23_GT00 = R20C23_GT00;
assign R17C23_GT10 = R20C23_GT10;
assign R18C23_GT00 = R20C23_GT00;
assign R18C23_GT10 = R20C23_GT10;
assign R21C23_GT00 = R20C23_GT00;
assign R21C23_GT10 = R20C23_GT10;
assign R22C23_GT00 = R20C23_GT00;
assign R22C23_GT10 = R20C23_GT10;
assign R23C23_GT00 = R20C23_GT00;
assign R23C23_GT10 = R20C23_GT10;
assign R24C23_GT00 = R20C23_GT00;
assign R24C23_GT10 = R20C23_GT10;
assign R25C23_GT00 = R20C23_GT00;
assign R25C23_GT10 = R20C23_GT10;
assign R26C23_GT00 = R20C23_GT00;
assign R26C23_GT10 = R20C23_GT10;
assign R27C23_GT00 = R20C23_GT00;
assign R27C23_GT10 = R20C23_GT10;
assign R11C24_GT00 = R20C24_GT00;
assign R11C24_GT10 = R20C24_GT10;
assign R12C24_GT00 = R20C24_GT00;
assign R12C24_GT10 = R20C24_GT10;
assign R13C24_GT00 = R20C24_GT00;
assign R13C24_GT10 = R20C24_GT10;
assign R14C24_GT00 = R20C24_GT00;
assign R14C24_GT10 = R20C24_GT10;
assign R15C24_GT00 = R20C24_GT00;
assign R15C24_GT10 = R20C24_GT10;
assign R16C24_GT00 = R20C24_GT00;
assign R16C24_GT10 = R20C24_GT10;
assign R17C24_GT00 = R20C24_GT00;
assign R17C24_GT10 = R20C24_GT10;
assign R18C24_GT00 = R20C24_GT00;
assign R18C24_GT10 = R20C24_GT10;
assign R21C24_GT00 = R20C24_GT00;
assign R21C24_GT10 = R20C24_GT10;
assign R22C24_GT00 = R20C24_GT00;
assign R22C24_GT10 = R20C24_GT10;
assign R23C24_GT00 = R20C24_GT00;
assign R23C24_GT10 = R20C24_GT10;
assign R24C24_GT00 = R20C24_GT00;
assign R24C24_GT10 = R20C24_GT10;
assign R25C24_GT00 = R20C24_GT00;
assign R25C24_GT10 = R20C24_GT10;
assign R26C24_GT00 = R20C24_GT00;
assign R26C24_GT10 = R20C24_GT10;
assign R27C24_GT00 = R20C24_GT00;
assign R27C24_GT10 = R20C24_GT10;
assign R11C25_GT00 = R20C25_GT00;
assign R11C25_GT10 = R20C25_GT10;
assign R12C25_GT00 = R20C25_GT00;
assign R12C25_GT10 = R20C25_GT10;
assign R13C25_GT00 = R20C25_GT00;
assign R13C25_GT10 = R20C25_GT10;
assign R14C25_GT00 = R20C25_GT00;
assign R14C25_GT10 = R20C25_GT10;
assign R15C25_GT00 = R20C25_GT00;
assign R15C25_GT10 = R20C25_GT10;
assign R16C25_GT00 = R20C25_GT00;
assign R16C25_GT10 = R20C25_GT10;
assign R17C25_GT00 = R20C25_GT00;
assign R17C25_GT10 = R20C25_GT10;
assign R18C25_GT00 = R20C25_GT00;
assign R18C25_GT10 = R20C25_GT10;
assign R21C25_GT00 = R20C25_GT00;
assign R21C25_GT10 = R20C25_GT10;
assign R22C25_GT00 = R20C25_GT00;
assign R22C25_GT10 = R20C25_GT10;
assign R23C25_GT00 = R20C25_GT00;
assign R23C25_GT10 = R20C25_GT10;
assign R24C25_GT00 = R20C25_GT00;
assign R24C25_GT10 = R20C25_GT10;
assign R25C25_GT00 = R20C25_GT00;
assign R25C25_GT10 = R20C25_GT10;
assign R26C25_GT00 = R20C25_GT00;
assign R26C25_GT10 = R20C25_GT10;
assign R27C25_GT00 = R20C25_GT00;
assign R27C25_GT10 = R20C25_GT10;
assign R11C26_GT00 = R20C26_GT00;
assign R11C26_GT10 = R20C26_GT10;
assign R12C26_GT00 = R20C26_GT00;
assign R12C26_GT10 = R20C26_GT10;
assign R13C26_GT00 = R20C26_GT00;
assign R13C26_GT10 = R20C26_GT10;
assign R14C26_GT00 = R20C26_GT00;
assign R14C26_GT10 = R20C26_GT10;
assign R15C26_GT00 = R20C26_GT00;
assign R15C26_GT10 = R20C26_GT10;
assign R16C26_GT00 = R20C26_GT00;
assign R16C26_GT10 = R20C26_GT10;
assign R17C26_GT00 = R20C26_GT00;
assign R17C26_GT10 = R20C26_GT10;
assign R18C26_GT00 = R20C26_GT00;
assign R18C26_GT10 = R20C26_GT10;
assign R21C26_GT00 = R20C26_GT00;
assign R21C26_GT10 = R20C26_GT10;
assign R22C26_GT00 = R20C26_GT00;
assign R22C26_GT10 = R20C26_GT10;
assign R23C26_GT00 = R20C26_GT00;
assign R23C26_GT10 = R20C26_GT10;
assign R24C26_GT00 = R20C26_GT00;
assign R24C26_GT10 = R20C26_GT10;
assign R25C26_GT00 = R20C26_GT00;
assign R25C26_GT10 = R20C26_GT10;
assign R26C26_GT00 = R20C26_GT00;
assign R26C26_GT10 = R20C26_GT10;
assign R27C26_GT00 = R20C26_GT00;
assign R27C26_GT10 = R20C26_GT10;
assign R11C27_GT00 = R20C27_GT00;
assign R11C27_GT10 = R20C27_GT10;
assign R12C27_GT00 = R20C27_GT00;
assign R12C27_GT10 = R20C27_GT10;
assign R13C27_GT00 = R20C27_GT00;
assign R13C27_GT10 = R20C27_GT10;
assign R14C27_GT00 = R20C27_GT00;
assign R14C27_GT10 = R20C27_GT10;
assign R15C27_GT00 = R20C27_GT00;
assign R15C27_GT10 = R20C27_GT10;
assign R16C27_GT00 = R20C27_GT00;
assign R16C27_GT10 = R20C27_GT10;
assign R17C27_GT00 = R20C27_GT00;
assign R17C27_GT10 = R20C27_GT10;
assign R18C27_GT00 = R20C27_GT00;
assign R18C27_GT10 = R20C27_GT10;
assign R21C27_GT00 = R20C27_GT00;
assign R21C27_GT10 = R20C27_GT10;
assign R22C27_GT00 = R20C27_GT00;
assign R22C27_GT10 = R20C27_GT10;
assign R23C27_GT00 = R20C27_GT00;
assign R23C27_GT10 = R20C27_GT10;
assign R24C27_GT00 = R20C27_GT00;
assign R24C27_GT10 = R20C27_GT10;
assign R25C27_GT00 = R20C27_GT00;
assign R25C27_GT10 = R20C27_GT10;
assign R26C27_GT00 = R20C27_GT00;
assign R26C27_GT10 = R20C27_GT10;
assign R27C27_GT00 = R20C27_GT00;
assign R27C27_GT10 = R20C27_GT10;
assign R11C28_GT00 = R20C28_GT00;
assign R11C28_GT10 = R20C28_GT10;
assign R12C28_GT00 = R20C28_GT00;
assign R12C28_GT10 = R20C28_GT10;
assign R13C28_GT00 = R20C28_GT00;
assign R13C28_GT10 = R20C28_GT10;
assign R14C28_GT00 = R20C28_GT00;
assign R14C28_GT10 = R20C28_GT10;
assign R15C28_GT00 = R20C28_GT00;
assign R15C28_GT10 = R20C28_GT10;
assign R16C28_GT00 = R20C28_GT00;
assign R16C28_GT10 = R20C28_GT10;
assign R17C28_GT00 = R20C28_GT00;
assign R17C28_GT10 = R20C28_GT10;
assign R18C28_GT00 = R20C28_GT00;
assign R18C28_GT10 = R20C28_GT10;
assign R21C28_GT00 = R20C28_GT00;
assign R21C28_GT10 = R20C28_GT10;
assign R22C28_GT00 = R20C28_GT00;
assign R22C28_GT10 = R20C28_GT10;
assign R23C28_GT00 = R20C28_GT00;
assign R23C28_GT10 = R20C28_GT10;
assign R24C28_GT00 = R20C28_GT00;
assign R24C28_GT10 = R20C28_GT10;
assign R25C28_GT00 = R20C28_GT00;
assign R25C28_GT10 = R20C28_GT10;
assign R26C28_GT00 = R20C28_GT00;
assign R26C28_GT10 = R20C28_GT10;
assign R27C28_GT00 = R20C28_GT00;
assign R27C28_GT10 = R20C28_GT10;
assign R3C33_GT00 = R2C33_GT00;
assign R3C33_GT10 = R2C33_GT10;
assign R4C33_GT00 = R2C33_GT00;
assign R4C33_GT10 = R2C33_GT10;
assign R5C33_GT00 = R2C33_GT00;
assign R5C33_GT10 = R2C33_GT10;
assign R6C33_GT00 = R2C33_GT00;
assign R6C33_GT10 = R2C33_GT10;
assign R7C33_GT00 = R2C33_GT00;
assign R7C33_GT10 = R2C33_GT10;
assign R8C33_GT00 = R2C33_GT00;
assign R8C33_GT10 = R2C33_GT10;
assign R9C33_GT00 = R2C33_GT00;
assign R9C33_GT10 = R2C33_GT10;
assign R3C34_GT00 = R2C34_GT00;
assign R3C34_GT10 = R2C34_GT10;
assign R4C34_GT00 = R2C34_GT00;
assign R4C34_GT10 = R2C34_GT10;
assign R5C34_GT00 = R2C34_GT00;
assign R5C34_GT10 = R2C34_GT10;
assign R6C34_GT00 = R2C34_GT00;
assign R6C34_GT10 = R2C34_GT10;
assign R7C34_GT00 = R2C34_GT00;
assign R7C34_GT10 = R2C34_GT10;
assign R8C34_GT00 = R2C34_GT00;
assign R8C34_GT10 = R2C34_GT10;
assign R9C34_GT00 = R2C34_GT00;
assign R9C34_GT10 = R2C34_GT10;
assign R3C35_GT00 = R2C35_GT00;
assign R3C35_GT10 = R2C35_GT10;
assign R4C35_GT00 = R2C35_GT00;
assign R4C35_GT10 = R2C35_GT10;
assign R5C35_GT00 = R2C35_GT00;
assign R5C35_GT10 = R2C35_GT10;
assign R6C35_GT00 = R2C35_GT00;
assign R6C35_GT10 = R2C35_GT10;
assign R7C35_GT00 = R2C35_GT00;
assign R7C35_GT10 = R2C35_GT10;
assign R8C35_GT00 = R2C35_GT00;
assign R8C35_GT10 = R2C35_GT10;
assign R9C35_GT00 = R2C35_GT00;
assign R9C35_GT10 = R2C35_GT10;
assign R3C36_GT00 = R2C36_GT00;
assign R3C36_GT10 = R2C36_GT10;
assign R4C36_GT00 = R2C36_GT00;
assign R4C36_GT10 = R2C36_GT10;
assign R5C36_GT00 = R2C36_GT00;
assign R5C36_GT10 = R2C36_GT10;
assign R6C36_GT00 = R2C36_GT00;
assign R6C36_GT10 = R2C36_GT10;
assign R7C36_GT00 = R2C36_GT00;
assign R7C36_GT10 = R2C36_GT10;
assign R8C36_GT00 = R2C36_GT00;
assign R8C36_GT10 = R2C36_GT10;
assign R9C36_GT00 = R2C36_GT00;
assign R9C36_GT10 = R2C36_GT10;
assign R3C37_GT00 = R2C37_GT00;
assign R3C37_GT10 = R2C37_GT10;
assign R4C37_GT00 = R2C37_GT00;
assign R4C37_GT10 = R2C37_GT10;
assign R5C37_GT00 = R2C37_GT00;
assign R5C37_GT10 = R2C37_GT10;
assign R6C37_GT00 = R2C37_GT00;
assign R6C37_GT10 = R2C37_GT10;
assign R7C37_GT00 = R2C37_GT00;
assign R7C37_GT10 = R2C37_GT10;
assign R8C37_GT00 = R2C37_GT00;
assign R8C37_GT10 = R2C37_GT10;
assign R9C37_GT00 = R2C37_GT00;
assign R9C37_GT10 = R2C37_GT10;
assign R3C38_GT00 = R2C38_GT00;
assign R3C38_GT10 = R2C38_GT10;
assign R4C38_GT00 = R2C38_GT00;
assign R4C38_GT10 = R2C38_GT10;
assign R5C38_GT00 = R2C38_GT00;
assign R5C38_GT10 = R2C38_GT10;
assign R6C38_GT00 = R2C38_GT00;
assign R6C38_GT10 = R2C38_GT10;
assign R7C38_GT00 = R2C38_GT00;
assign R7C38_GT10 = R2C38_GT10;
assign R8C38_GT00 = R2C38_GT00;
assign R8C38_GT10 = R2C38_GT10;
assign R9C38_GT00 = R2C38_GT00;
assign R9C38_GT10 = R2C38_GT10;
assign R3C39_GT00 = R2C39_GT00;
assign R3C39_GT10 = R2C39_GT10;
assign R4C39_GT00 = R2C39_GT00;
assign R4C39_GT10 = R2C39_GT10;
assign R5C39_GT00 = R2C39_GT00;
assign R5C39_GT10 = R2C39_GT10;
assign R6C39_GT00 = R2C39_GT00;
assign R6C39_GT10 = R2C39_GT10;
assign R7C39_GT00 = R2C39_GT00;
assign R7C39_GT10 = R2C39_GT10;
assign R8C39_GT00 = R2C39_GT00;
assign R8C39_GT10 = R2C39_GT10;
assign R9C39_GT00 = R2C39_GT00;
assign R9C39_GT10 = R2C39_GT10;
assign R3C40_GT00 = R2C40_GT00;
assign R3C40_GT10 = R2C40_GT10;
assign R4C40_GT00 = R2C40_GT00;
assign R4C40_GT10 = R2C40_GT10;
assign R5C40_GT00 = R2C40_GT00;
assign R5C40_GT10 = R2C40_GT10;
assign R6C40_GT00 = R2C40_GT00;
assign R6C40_GT10 = R2C40_GT10;
assign R7C40_GT00 = R2C40_GT00;
assign R7C40_GT10 = R2C40_GT10;
assign R8C40_GT00 = R2C40_GT00;
assign R8C40_GT10 = R2C40_GT10;
assign R9C40_GT00 = R2C40_GT00;
assign R9C40_GT10 = R2C40_GT10;
assign R3C41_GT00 = R2C41_GT00;
assign R3C41_GT10 = R2C41_GT10;
assign R4C41_GT00 = R2C41_GT00;
assign R4C41_GT10 = R2C41_GT10;
assign R5C41_GT00 = R2C41_GT00;
assign R5C41_GT10 = R2C41_GT10;
assign R6C41_GT00 = R2C41_GT00;
assign R6C41_GT10 = R2C41_GT10;
assign R7C41_GT00 = R2C41_GT00;
assign R7C41_GT10 = R2C41_GT10;
assign R8C41_GT00 = R2C41_GT00;
assign R8C41_GT10 = R2C41_GT10;
assign R9C41_GT00 = R2C41_GT00;
assign R9C41_GT10 = R2C41_GT10;
assign R3C42_GT00 = R2C42_GT00;
assign R3C42_GT10 = R2C42_GT10;
assign R4C42_GT00 = R2C42_GT00;
assign R4C42_GT10 = R2C42_GT10;
assign R5C42_GT00 = R2C42_GT00;
assign R5C42_GT10 = R2C42_GT10;
assign R6C42_GT00 = R2C42_GT00;
assign R6C42_GT10 = R2C42_GT10;
assign R7C42_GT00 = R2C42_GT00;
assign R7C42_GT10 = R2C42_GT10;
assign R8C42_GT00 = R2C42_GT00;
assign R8C42_GT10 = R2C42_GT10;
assign R9C42_GT00 = R2C42_GT00;
assign R9C42_GT10 = R2C42_GT10;
assign R3C43_GT00 = R2C43_GT00;
assign R3C43_GT10 = R2C43_GT10;
assign R4C43_GT00 = R2C43_GT00;
assign R4C43_GT10 = R2C43_GT10;
assign R5C43_GT00 = R2C43_GT00;
assign R5C43_GT10 = R2C43_GT10;
assign R6C43_GT00 = R2C43_GT00;
assign R6C43_GT10 = R2C43_GT10;
assign R7C43_GT00 = R2C43_GT00;
assign R7C43_GT10 = R2C43_GT10;
assign R8C43_GT00 = R2C43_GT00;
assign R8C43_GT10 = R2C43_GT10;
assign R9C43_GT00 = R2C43_GT00;
assign R9C43_GT10 = R2C43_GT10;
assign R3C44_GT00 = R2C44_GT00;
assign R3C44_GT10 = R2C44_GT10;
assign R4C44_GT00 = R2C44_GT00;
assign R4C44_GT10 = R2C44_GT10;
assign R5C44_GT00 = R2C44_GT00;
assign R5C44_GT10 = R2C44_GT10;
assign R6C44_GT00 = R2C44_GT00;
assign R6C44_GT10 = R2C44_GT10;
assign R7C44_GT00 = R2C44_GT00;
assign R7C44_GT10 = R2C44_GT10;
assign R8C44_GT00 = R2C44_GT00;
assign R8C44_GT10 = R2C44_GT10;
assign R9C44_GT00 = R2C44_GT00;
assign R9C44_GT10 = R2C44_GT10;
assign R3C45_GT00 = R2C45_GT00;
assign R3C45_GT10 = R2C45_GT10;
assign R4C45_GT00 = R2C45_GT00;
assign R4C45_GT10 = R2C45_GT10;
assign R5C45_GT00 = R2C45_GT00;
assign R5C45_GT10 = R2C45_GT10;
assign R6C45_GT00 = R2C45_GT00;
assign R6C45_GT10 = R2C45_GT10;
assign R7C45_GT00 = R2C45_GT00;
assign R7C45_GT10 = R2C45_GT10;
assign R8C45_GT00 = R2C45_GT00;
assign R8C45_GT10 = R2C45_GT10;
assign R9C45_GT00 = R2C45_GT00;
assign R9C45_GT10 = R2C45_GT10;
assign R3C46_GT00 = R2C46_GT00;
assign R3C46_GT10 = R2C46_GT10;
assign R4C46_GT00 = R2C46_GT00;
assign R4C46_GT10 = R2C46_GT10;
assign R5C46_GT00 = R2C46_GT00;
assign R5C46_GT10 = R2C46_GT10;
assign R6C46_GT00 = R2C46_GT00;
assign R6C46_GT10 = R2C46_GT10;
assign R7C46_GT00 = R2C46_GT00;
assign R7C46_GT10 = R2C46_GT10;
assign R8C46_GT00 = R2C46_GT00;
assign R8C46_GT10 = R2C46_GT10;
assign R9C46_GT00 = R2C46_GT00;
assign R9C46_GT10 = R2C46_GT10;
assign R3C29_GT00 = R2C29_GT00;
assign R3C29_GT10 = R2C29_GT10;
assign R4C29_GT00 = R2C29_GT00;
assign R4C29_GT10 = R2C29_GT10;
assign R5C29_GT00 = R2C29_GT00;
assign R5C29_GT10 = R2C29_GT10;
assign R6C29_GT00 = R2C29_GT00;
assign R6C29_GT10 = R2C29_GT10;
assign R7C29_GT00 = R2C29_GT00;
assign R7C29_GT10 = R2C29_GT10;
assign R8C29_GT00 = R2C29_GT00;
assign R8C29_GT10 = R2C29_GT10;
assign R9C29_GT00 = R2C29_GT00;
assign R9C29_GT10 = R2C29_GT10;
assign R3C30_GT00 = R2C30_GT00;
assign R3C30_GT10 = R2C30_GT10;
assign R4C30_GT00 = R2C30_GT00;
assign R4C30_GT10 = R2C30_GT10;
assign R5C30_GT00 = R2C30_GT00;
assign R5C30_GT10 = R2C30_GT10;
assign R6C30_GT00 = R2C30_GT00;
assign R6C30_GT10 = R2C30_GT10;
assign R7C30_GT00 = R2C30_GT00;
assign R7C30_GT10 = R2C30_GT10;
assign R8C30_GT00 = R2C30_GT00;
assign R8C30_GT10 = R2C30_GT10;
assign R9C30_GT00 = R2C30_GT00;
assign R9C30_GT10 = R2C30_GT10;
assign R3C31_GT00 = R2C31_GT00;
assign R3C31_GT10 = R2C31_GT10;
assign R4C31_GT00 = R2C31_GT00;
assign R4C31_GT10 = R2C31_GT10;
assign R5C31_GT00 = R2C31_GT00;
assign R5C31_GT10 = R2C31_GT10;
assign R6C31_GT00 = R2C31_GT00;
assign R6C31_GT10 = R2C31_GT10;
assign R7C31_GT00 = R2C31_GT00;
assign R7C31_GT10 = R2C31_GT10;
assign R8C31_GT00 = R2C31_GT00;
assign R8C31_GT10 = R2C31_GT10;
assign R9C31_GT00 = R2C31_GT00;
assign R9C31_GT10 = R2C31_GT10;
assign R3C32_GT00 = R2C32_GT00;
assign R3C32_GT10 = R2C32_GT10;
assign R4C32_GT00 = R2C32_GT00;
assign R4C32_GT10 = R2C32_GT10;
assign R5C32_GT00 = R2C32_GT00;
assign R5C32_GT10 = R2C32_GT10;
assign R6C32_GT00 = R2C32_GT00;
assign R6C32_GT10 = R2C32_GT10;
assign R7C32_GT00 = R2C32_GT00;
assign R7C32_GT10 = R2C32_GT10;
assign R8C32_GT00 = R2C32_GT00;
assign R8C32_GT10 = R2C32_GT10;
assign R9C32_GT00 = R2C32_GT00;
assign R9C32_GT10 = R2C32_GT10;
assign R11C33_GT00 = R20C33_GT00;
assign R11C33_GT10 = R20C33_GT10;
assign R12C33_GT00 = R20C33_GT00;
assign R12C33_GT10 = R20C33_GT10;
assign R13C33_GT00 = R20C33_GT00;
assign R13C33_GT10 = R20C33_GT10;
assign R14C33_GT00 = R20C33_GT00;
assign R14C33_GT10 = R20C33_GT10;
assign R15C33_GT00 = R20C33_GT00;
assign R15C33_GT10 = R20C33_GT10;
assign R16C33_GT00 = R20C33_GT00;
assign R16C33_GT10 = R20C33_GT10;
assign R17C33_GT00 = R20C33_GT00;
assign R17C33_GT10 = R20C33_GT10;
assign R18C33_GT00 = R20C33_GT00;
assign R18C33_GT10 = R20C33_GT10;
assign R21C33_GT00 = R20C33_GT00;
assign R21C33_GT10 = R20C33_GT10;
assign R22C33_GT00 = R20C33_GT00;
assign R22C33_GT10 = R20C33_GT10;
assign R23C33_GT00 = R20C33_GT00;
assign R23C33_GT10 = R20C33_GT10;
assign R24C33_GT00 = R20C33_GT00;
assign R24C33_GT10 = R20C33_GT10;
assign R25C33_GT00 = R20C33_GT00;
assign R25C33_GT10 = R20C33_GT10;
assign R26C33_GT00 = R20C33_GT00;
assign R26C33_GT10 = R20C33_GT10;
assign R27C33_GT00 = R20C33_GT00;
assign R27C33_GT10 = R20C33_GT10;
assign R11C34_GT00 = R20C34_GT00;
assign R11C34_GT10 = R20C34_GT10;
assign R12C34_GT00 = R20C34_GT00;
assign R12C34_GT10 = R20C34_GT10;
assign R13C34_GT00 = R20C34_GT00;
assign R13C34_GT10 = R20C34_GT10;
assign R14C34_GT00 = R20C34_GT00;
assign R14C34_GT10 = R20C34_GT10;
assign R15C34_GT00 = R20C34_GT00;
assign R15C34_GT10 = R20C34_GT10;
assign R16C34_GT00 = R20C34_GT00;
assign R16C34_GT10 = R20C34_GT10;
assign R17C34_GT00 = R20C34_GT00;
assign R17C34_GT10 = R20C34_GT10;
assign R18C34_GT00 = R20C34_GT00;
assign R18C34_GT10 = R20C34_GT10;
assign R21C34_GT00 = R20C34_GT00;
assign R21C34_GT10 = R20C34_GT10;
assign R22C34_GT00 = R20C34_GT00;
assign R22C34_GT10 = R20C34_GT10;
assign R23C34_GT00 = R20C34_GT00;
assign R23C34_GT10 = R20C34_GT10;
assign R24C34_GT00 = R20C34_GT00;
assign R24C34_GT10 = R20C34_GT10;
assign R25C34_GT00 = R20C34_GT00;
assign R25C34_GT10 = R20C34_GT10;
assign R26C34_GT00 = R20C34_GT00;
assign R26C34_GT10 = R20C34_GT10;
assign R27C34_GT00 = R20C34_GT00;
assign R27C34_GT10 = R20C34_GT10;
assign R11C35_GT00 = R20C35_GT00;
assign R11C35_GT10 = R20C35_GT10;
assign R12C35_GT00 = R20C35_GT00;
assign R12C35_GT10 = R20C35_GT10;
assign R13C35_GT00 = R20C35_GT00;
assign R13C35_GT10 = R20C35_GT10;
assign R14C35_GT00 = R20C35_GT00;
assign R14C35_GT10 = R20C35_GT10;
assign R15C35_GT00 = R20C35_GT00;
assign R15C35_GT10 = R20C35_GT10;
assign R16C35_GT00 = R20C35_GT00;
assign R16C35_GT10 = R20C35_GT10;
assign R17C35_GT00 = R20C35_GT00;
assign R17C35_GT10 = R20C35_GT10;
assign R18C35_GT00 = R20C35_GT00;
assign R18C35_GT10 = R20C35_GT10;
assign R21C35_GT00 = R20C35_GT00;
assign R21C35_GT10 = R20C35_GT10;
assign R22C35_GT00 = R20C35_GT00;
assign R22C35_GT10 = R20C35_GT10;
assign R23C35_GT00 = R20C35_GT00;
assign R23C35_GT10 = R20C35_GT10;
assign R24C35_GT00 = R20C35_GT00;
assign R24C35_GT10 = R20C35_GT10;
assign R25C35_GT00 = R20C35_GT00;
assign R25C35_GT10 = R20C35_GT10;
assign R26C35_GT00 = R20C35_GT00;
assign R26C35_GT10 = R20C35_GT10;
assign R27C35_GT00 = R20C35_GT00;
assign R27C35_GT10 = R20C35_GT10;
assign R11C36_GT00 = R20C36_GT00;
assign R11C36_GT10 = R20C36_GT10;
assign R12C36_GT00 = R20C36_GT00;
assign R12C36_GT10 = R20C36_GT10;
assign R13C36_GT00 = R20C36_GT00;
assign R13C36_GT10 = R20C36_GT10;
assign R14C36_GT00 = R20C36_GT00;
assign R14C36_GT10 = R20C36_GT10;
assign R15C36_GT00 = R20C36_GT00;
assign R15C36_GT10 = R20C36_GT10;
assign R16C36_GT00 = R20C36_GT00;
assign R16C36_GT10 = R20C36_GT10;
assign R17C36_GT00 = R20C36_GT00;
assign R17C36_GT10 = R20C36_GT10;
assign R18C36_GT00 = R20C36_GT00;
assign R18C36_GT10 = R20C36_GT10;
assign R21C36_GT00 = R20C36_GT00;
assign R21C36_GT10 = R20C36_GT10;
assign R22C36_GT00 = R20C36_GT00;
assign R22C36_GT10 = R20C36_GT10;
assign R23C36_GT00 = R20C36_GT00;
assign R23C36_GT10 = R20C36_GT10;
assign R24C36_GT00 = R20C36_GT00;
assign R24C36_GT10 = R20C36_GT10;
assign R25C36_GT00 = R20C36_GT00;
assign R25C36_GT10 = R20C36_GT10;
assign R26C36_GT00 = R20C36_GT00;
assign R26C36_GT10 = R20C36_GT10;
assign R27C36_GT00 = R20C36_GT00;
assign R27C36_GT10 = R20C36_GT10;
assign R11C37_GT00 = R20C37_GT00;
assign R11C37_GT10 = R20C37_GT10;
assign R12C37_GT00 = R20C37_GT00;
assign R12C37_GT10 = R20C37_GT10;
assign R13C37_GT00 = R20C37_GT00;
assign R13C37_GT10 = R20C37_GT10;
assign R14C37_GT00 = R20C37_GT00;
assign R14C37_GT10 = R20C37_GT10;
assign R15C37_GT00 = R20C37_GT00;
assign R15C37_GT10 = R20C37_GT10;
assign R16C37_GT00 = R20C37_GT00;
assign R16C37_GT10 = R20C37_GT10;
assign R17C37_GT00 = R20C37_GT00;
assign R17C37_GT10 = R20C37_GT10;
assign R18C37_GT00 = R20C37_GT00;
assign R18C37_GT10 = R20C37_GT10;
assign R21C37_GT00 = R20C37_GT00;
assign R21C37_GT10 = R20C37_GT10;
assign R22C37_GT00 = R20C37_GT00;
assign R22C37_GT10 = R20C37_GT10;
assign R23C37_GT00 = R20C37_GT00;
assign R23C37_GT10 = R20C37_GT10;
assign R24C37_GT00 = R20C37_GT00;
assign R24C37_GT10 = R20C37_GT10;
assign R25C37_GT00 = R20C37_GT00;
assign R25C37_GT10 = R20C37_GT10;
assign R26C37_GT00 = R20C37_GT00;
assign R26C37_GT10 = R20C37_GT10;
assign R27C37_GT00 = R20C37_GT00;
assign R27C37_GT10 = R20C37_GT10;
assign R11C38_GT00 = R20C38_GT00;
assign R11C38_GT10 = R20C38_GT10;
assign R12C38_GT00 = R20C38_GT00;
assign R12C38_GT10 = R20C38_GT10;
assign R13C38_GT00 = R20C38_GT00;
assign R13C38_GT10 = R20C38_GT10;
assign R14C38_GT00 = R20C38_GT00;
assign R14C38_GT10 = R20C38_GT10;
assign R15C38_GT00 = R20C38_GT00;
assign R15C38_GT10 = R20C38_GT10;
assign R16C38_GT00 = R20C38_GT00;
assign R16C38_GT10 = R20C38_GT10;
assign R17C38_GT00 = R20C38_GT00;
assign R17C38_GT10 = R20C38_GT10;
assign R18C38_GT00 = R20C38_GT00;
assign R18C38_GT10 = R20C38_GT10;
assign R21C38_GT00 = R20C38_GT00;
assign R21C38_GT10 = R20C38_GT10;
assign R22C38_GT00 = R20C38_GT00;
assign R22C38_GT10 = R20C38_GT10;
assign R23C38_GT00 = R20C38_GT00;
assign R23C38_GT10 = R20C38_GT10;
assign R24C38_GT00 = R20C38_GT00;
assign R24C38_GT10 = R20C38_GT10;
assign R25C38_GT00 = R20C38_GT00;
assign R25C38_GT10 = R20C38_GT10;
assign R26C38_GT00 = R20C38_GT00;
assign R26C38_GT10 = R20C38_GT10;
assign R27C38_GT00 = R20C38_GT00;
assign R27C38_GT10 = R20C38_GT10;
assign R11C39_GT00 = R20C39_GT00;
assign R11C39_GT10 = R20C39_GT10;
assign R12C39_GT00 = R20C39_GT00;
assign R12C39_GT10 = R20C39_GT10;
assign R13C39_GT00 = R20C39_GT00;
assign R13C39_GT10 = R20C39_GT10;
assign R14C39_GT00 = R20C39_GT00;
assign R14C39_GT10 = R20C39_GT10;
assign R15C39_GT00 = R20C39_GT00;
assign R15C39_GT10 = R20C39_GT10;
assign R16C39_GT00 = R20C39_GT00;
assign R16C39_GT10 = R20C39_GT10;
assign R17C39_GT00 = R20C39_GT00;
assign R17C39_GT10 = R20C39_GT10;
assign R18C39_GT00 = R20C39_GT00;
assign R18C39_GT10 = R20C39_GT10;
assign R21C39_GT00 = R20C39_GT00;
assign R21C39_GT10 = R20C39_GT10;
assign R22C39_GT00 = R20C39_GT00;
assign R22C39_GT10 = R20C39_GT10;
assign R23C39_GT00 = R20C39_GT00;
assign R23C39_GT10 = R20C39_GT10;
assign R24C39_GT00 = R20C39_GT00;
assign R24C39_GT10 = R20C39_GT10;
assign R25C39_GT00 = R20C39_GT00;
assign R25C39_GT10 = R20C39_GT10;
assign R26C39_GT00 = R20C39_GT00;
assign R26C39_GT10 = R20C39_GT10;
assign R27C39_GT00 = R20C39_GT00;
assign R27C39_GT10 = R20C39_GT10;
assign R11C40_GT00 = R20C40_GT00;
assign R11C40_GT10 = R20C40_GT10;
assign R12C40_GT00 = R20C40_GT00;
assign R12C40_GT10 = R20C40_GT10;
assign R13C40_GT00 = R20C40_GT00;
assign R13C40_GT10 = R20C40_GT10;
assign R14C40_GT00 = R20C40_GT00;
assign R14C40_GT10 = R20C40_GT10;
assign R15C40_GT00 = R20C40_GT00;
assign R15C40_GT10 = R20C40_GT10;
assign R16C40_GT00 = R20C40_GT00;
assign R16C40_GT10 = R20C40_GT10;
assign R17C40_GT00 = R20C40_GT00;
assign R17C40_GT10 = R20C40_GT10;
assign R18C40_GT00 = R20C40_GT00;
assign R18C40_GT10 = R20C40_GT10;
assign R21C40_GT00 = R20C40_GT00;
assign R21C40_GT10 = R20C40_GT10;
assign R22C40_GT00 = R20C40_GT00;
assign R22C40_GT10 = R20C40_GT10;
assign R23C40_GT00 = R20C40_GT00;
assign R23C40_GT10 = R20C40_GT10;
assign R24C40_GT00 = R20C40_GT00;
assign R24C40_GT10 = R20C40_GT10;
assign R25C40_GT00 = R20C40_GT00;
assign R25C40_GT10 = R20C40_GT10;
assign R26C40_GT00 = R20C40_GT00;
assign R26C40_GT10 = R20C40_GT10;
assign R27C40_GT00 = R20C40_GT00;
assign R27C40_GT10 = R20C40_GT10;
assign R11C41_GT00 = R20C41_GT00;
assign R11C41_GT10 = R20C41_GT10;
assign R12C41_GT00 = R20C41_GT00;
assign R12C41_GT10 = R20C41_GT10;
assign R13C41_GT00 = R20C41_GT00;
assign R13C41_GT10 = R20C41_GT10;
assign R14C41_GT00 = R20C41_GT00;
assign R14C41_GT10 = R20C41_GT10;
assign R15C41_GT00 = R20C41_GT00;
assign R15C41_GT10 = R20C41_GT10;
assign R16C41_GT00 = R20C41_GT00;
assign R16C41_GT10 = R20C41_GT10;
assign R17C41_GT00 = R20C41_GT00;
assign R17C41_GT10 = R20C41_GT10;
assign R18C41_GT00 = R20C41_GT00;
assign R18C41_GT10 = R20C41_GT10;
assign R21C41_GT00 = R20C41_GT00;
assign R21C41_GT10 = R20C41_GT10;
assign R22C41_GT00 = R20C41_GT00;
assign R22C41_GT10 = R20C41_GT10;
assign R23C41_GT00 = R20C41_GT00;
assign R23C41_GT10 = R20C41_GT10;
assign R24C41_GT00 = R20C41_GT00;
assign R24C41_GT10 = R20C41_GT10;
assign R25C41_GT00 = R20C41_GT00;
assign R25C41_GT10 = R20C41_GT10;
assign R26C41_GT00 = R20C41_GT00;
assign R26C41_GT10 = R20C41_GT10;
assign R27C41_GT00 = R20C41_GT00;
assign R27C41_GT10 = R20C41_GT10;
assign R11C42_GT00 = R20C42_GT00;
assign R11C42_GT10 = R20C42_GT10;
assign R12C42_GT00 = R20C42_GT00;
assign R12C42_GT10 = R20C42_GT10;
assign R13C42_GT00 = R20C42_GT00;
assign R13C42_GT10 = R20C42_GT10;
assign R14C42_GT00 = R20C42_GT00;
assign R14C42_GT10 = R20C42_GT10;
assign R15C42_GT00 = R20C42_GT00;
assign R15C42_GT10 = R20C42_GT10;
assign R16C42_GT00 = R20C42_GT00;
assign R16C42_GT10 = R20C42_GT10;
assign R17C42_GT00 = R20C42_GT00;
assign R17C42_GT10 = R20C42_GT10;
assign R18C42_GT00 = R20C42_GT00;
assign R18C42_GT10 = R20C42_GT10;
assign R21C42_GT00 = R20C42_GT00;
assign R21C42_GT10 = R20C42_GT10;
assign R22C42_GT00 = R20C42_GT00;
assign R22C42_GT10 = R20C42_GT10;
assign R23C42_GT00 = R20C42_GT00;
assign R23C42_GT10 = R20C42_GT10;
assign R24C42_GT00 = R20C42_GT00;
assign R24C42_GT10 = R20C42_GT10;
assign R25C42_GT00 = R20C42_GT00;
assign R25C42_GT10 = R20C42_GT10;
assign R26C42_GT00 = R20C42_GT00;
assign R26C42_GT10 = R20C42_GT10;
assign R27C42_GT00 = R20C42_GT00;
assign R27C42_GT10 = R20C42_GT10;
assign R11C43_GT00 = R20C43_GT00;
assign R11C43_GT10 = R20C43_GT10;
assign R12C43_GT00 = R20C43_GT00;
assign R12C43_GT10 = R20C43_GT10;
assign R13C43_GT00 = R20C43_GT00;
assign R13C43_GT10 = R20C43_GT10;
assign R14C43_GT00 = R20C43_GT00;
assign R14C43_GT10 = R20C43_GT10;
assign R15C43_GT00 = R20C43_GT00;
assign R15C43_GT10 = R20C43_GT10;
assign R16C43_GT00 = R20C43_GT00;
assign R16C43_GT10 = R20C43_GT10;
assign R17C43_GT00 = R20C43_GT00;
assign R17C43_GT10 = R20C43_GT10;
assign R18C43_GT00 = R20C43_GT00;
assign R18C43_GT10 = R20C43_GT10;
assign R21C43_GT00 = R20C43_GT00;
assign R21C43_GT10 = R20C43_GT10;
assign R22C43_GT00 = R20C43_GT00;
assign R22C43_GT10 = R20C43_GT10;
assign R23C43_GT00 = R20C43_GT00;
assign R23C43_GT10 = R20C43_GT10;
assign R24C43_GT00 = R20C43_GT00;
assign R24C43_GT10 = R20C43_GT10;
assign R25C43_GT00 = R20C43_GT00;
assign R25C43_GT10 = R20C43_GT10;
assign R26C43_GT00 = R20C43_GT00;
assign R26C43_GT10 = R20C43_GT10;
assign R27C43_GT00 = R20C43_GT00;
assign R27C43_GT10 = R20C43_GT10;
assign R11C44_GT00 = R20C44_GT00;
assign R11C44_GT10 = R20C44_GT10;
assign R12C44_GT00 = R20C44_GT00;
assign R12C44_GT10 = R20C44_GT10;
assign R13C44_GT00 = R20C44_GT00;
assign R13C44_GT10 = R20C44_GT10;
assign R14C44_GT00 = R20C44_GT00;
assign R14C44_GT10 = R20C44_GT10;
assign R15C44_GT00 = R20C44_GT00;
assign R15C44_GT10 = R20C44_GT10;
assign R16C44_GT00 = R20C44_GT00;
assign R16C44_GT10 = R20C44_GT10;
assign R17C44_GT00 = R20C44_GT00;
assign R17C44_GT10 = R20C44_GT10;
assign R18C44_GT00 = R20C44_GT00;
assign R18C44_GT10 = R20C44_GT10;
assign R21C44_GT00 = R20C44_GT00;
assign R21C44_GT10 = R20C44_GT10;
assign R22C44_GT00 = R20C44_GT00;
assign R22C44_GT10 = R20C44_GT10;
assign R23C44_GT00 = R20C44_GT00;
assign R23C44_GT10 = R20C44_GT10;
assign R24C44_GT00 = R20C44_GT00;
assign R24C44_GT10 = R20C44_GT10;
assign R25C44_GT00 = R20C44_GT00;
assign R25C44_GT10 = R20C44_GT10;
assign R26C44_GT00 = R20C44_GT00;
assign R26C44_GT10 = R20C44_GT10;
assign R27C44_GT00 = R20C44_GT00;
assign R27C44_GT10 = R20C44_GT10;
assign R11C45_GT00 = R20C45_GT00;
assign R11C45_GT10 = R20C45_GT10;
assign R12C45_GT00 = R20C45_GT00;
assign R12C45_GT10 = R20C45_GT10;
assign R13C45_GT00 = R20C45_GT00;
assign R13C45_GT10 = R20C45_GT10;
assign R14C45_GT00 = R20C45_GT00;
assign R14C45_GT10 = R20C45_GT10;
assign R15C45_GT00 = R20C45_GT00;
assign R15C45_GT10 = R20C45_GT10;
assign R16C45_GT00 = R20C45_GT00;
assign R16C45_GT10 = R20C45_GT10;
assign R17C45_GT00 = R20C45_GT00;
assign R17C45_GT10 = R20C45_GT10;
assign R18C45_GT00 = R20C45_GT00;
assign R18C45_GT10 = R20C45_GT10;
assign R21C45_GT00 = R20C45_GT00;
assign R21C45_GT10 = R20C45_GT10;
assign R22C45_GT00 = R20C45_GT00;
assign R22C45_GT10 = R20C45_GT10;
assign R23C45_GT00 = R20C45_GT00;
assign R23C45_GT10 = R20C45_GT10;
assign R24C45_GT00 = R20C45_GT00;
assign R24C45_GT10 = R20C45_GT10;
assign R25C45_GT00 = R20C45_GT00;
assign R25C45_GT10 = R20C45_GT10;
assign R26C45_GT00 = R20C45_GT00;
assign R26C45_GT10 = R20C45_GT10;
assign R27C45_GT00 = R20C45_GT00;
assign R27C45_GT10 = R20C45_GT10;
assign R11C46_GT00 = R20C46_GT00;
assign R11C46_GT10 = R20C46_GT10;
assign R12C46_GT00 = R20C46_GT00;
assign R12C46_GT10 = R20C46_GT10;
assign R13C46_GT00 = R20C46_GT00;
assign R13C46_GT10 = R20C46_GT10;
assign R14C46_GT00 = R20C46_GT00;
assign R14C46_GT10 = R20C46_GT10;
assign R15C46_GT00 = R20C46_GT00;
assign R15C46_GT10 = R20C46_GT10;
assign R16C46_GT00 = R20C46_GT00;
assign R16C46_GT10 = R20C46_GT10;
assign R17C46_GT00 = R20C46_GT00;
assign R17C46_GT10 = R20C46_GT10;
assign R18C46_GT00 = R20C46_GT00;
assign R18C46_GT10 = R20C46_GT10;
assign R21C46_GT00 = R20C46_GT00;
assign R21C46_GT10 = R20C46_GT10;
assign R22C46_GT00 = R20C46_GT00;
assign R22C46_GT10 = R20C46_GT10;
assign R23C46_GT00 = R20C46_GT00;
assign R23C46_GT10 = R20C46_GT10;
assign R24C46_GT00 = R20C46_GT00;
assign R24C46_GT10 = R20C46_GT10;
assign R25C46_GT00 = R20C46_GT00;
assign R25C46_GT10 = R20C46_GT10;
assign R26C46_GT00 = R20C46_GT00;
assign R26C46_GT10 = R20C46_GT10;
assign R27C46_GT00 = R20C46_GT00;
assign R27C46_GT10 = R20C46_GT10;
assign R11C29_GT00 = R20C29_GT00;
assign R11C29_GT10 = R20C29_GT10;
assign R12C29_GT00 = R20C29_GT00;
assign R12C29_GT10 = R20C29_GT10;
assign R13C29_GT00 = R20C29_GT00;
assign R13C29_GT10 = R20C29_GT10;
assign R14C29_GT00 = R20C29_GT00;
assign R14C29_GT10 = R20C29_GT10;
assign R15C29_GT00 = R20C29_GT00;
assign R15C29_GT10 = R20C29_GT10;
assign R16C29_GT00 = R20C29_GT00;
assign R16C29_GT10 = R20C29_GT10;
assign R17C29_GT00 = R20C29_GT00;
assign R17C29_GT10 = R20C29_GT10;
assign R18C29_GT00 = R20C29_GT00;
assign R18C29_GT10 = R20C29_GT10;
assign R21C29_GT00 = R20C29_GT00;
assign R21C29_GT10 = R20C29_GT10;
assign R22C29_GT00 = R20C29_GT00;
assign R22C29_GT10 = R20C29_GT10;
assign R23C29_GT00 = R20C29_GT00;
assign R23C29_GT10 = R20C29_GT10;
assign R24C29_GT00 = R20C29_GT00;
assign R24C29_GT10 = R20C29_GT10;
assign R25C29_GT00 = R20C29_GT00;
assign R25C29_GT10 = R20C29_GT10;
assign R26C29_GT00 = R20C29_GT00;
assign R26C29_GT10 = R20C29_GT10;
assign R27C29_GT00 = R20C29_GT00;
assign R27C29_GT10 = R20C29_GT10;
assign R11C30_GT00 = R20C30_GT00;
assign R11C30_GT10 = R20C30_GT10;
assign R12C30_GT00 = R20C30_GT00;
assign R12C30_GT10 = R20C30_GT10;
assign R13C30_GT00 = R20C30_GT00;
assign R13C30_GT10 = R20C30_GT10;
assign R14C30_GT00 = R20C30_GT00;
assign R14C30_GT10 = R20C30_GT10;
assign R15C30_GT00 = R20C30_GT00;
assign R15C30_GT10 = R20C30_GT10;
assign R16C30_GT00 = R20C30_GT00;
assign R16C30_GT10 = R20C30_GT10;
assign R17C30_GT00 = R20C30_GT00;
assign R17C30_GT10 = R20C30_GT10;
assign R18C30_GT00 = R20C30_GT00;
assign R18C30_GT10 = R20C30_GT10;
assign R21C30_GT00 = R20C30_GT00;
assign R21C30_GT10 = R20C30_GT10;
assign R22C30_GT00 = R20C30_GT00;
assign R22C30_GT10 = R20C30_GT10;
assign R23C30_GT00 = R20C30_GT00;
assign R23C30_GT10 = R20C30_GT10;
assign R24C30_GT00 = R20C30_GT00;
assign R24C30_GT10 = R20C30_GT10;
assign R25C30_GT00 = R20C30_GT00;
assign R25C30_GT10 = R20C30_GT10;
assign R26C30_GT00 = R20C30_GT00;
assign R26C30_GT10 = R20C30_GT10;
assign R27C30_GT00 = R20C30_GT00;
assign R27C30_GT10 = R20C30_GT10;
assign R11C31_GT00 = R20C31_GT00;
assign R11C31_GT10 = R20C31_GT10;
assign R12C31_GT00 = R20C31_GT00;
assign R12C31_GT10 = R20C31_GT10;
assign R13C31_GT00 = R20C31_GT00;
assign R13C31_GT10 = R20C31_GT10;
assign R14C31_GT00 = R20C31_GT00;
assign R14C31_GT10 = R20C31_GT10;
assign R15C31_GT00 = R20C31_GT00;
assign R15C31_GT10 = R20C31_GT10;
assign R16C31_GT00 = R20C31_GT00;
assign R16C31_GT10 = R20C31_GT10;
assign R17C31_GT00 = R20C31_GT00;
assign R17C31_GT10 = R20C31_GT10;
assign R18C31_GT00 = R20C31_GT00;
assign R18C31_GT10 = R20C31_GT10;
assign R21C31_GT00 = R20C31_GT00;
assign R21C31_GT10 = R20C31_GT10;
assign R22C31_GT00 = R20C31_GT00;
assign R22C31_GT10 = R20C31_GT10;
assign R23C31_GT00 = R20C31_GT00;
assign R23C31_GT10 = R20C31_GT10;
assign R24C31_GT00 = R20C31_GT00;
assign R24C31_GT10 = R20C31_GT10;
assign R25C31_GT00 = R20C31_GT00;
assign R25C31_GT10 = R20C31_GT10;
assign R26C31_GT00 = R20C31_GT00;
assign R26C31_GT10 = R20C31_GT10;
assign R27C31_GT00 = R20C31_GT00;
assign R27C31_GT10 = R20C31_GT10;
assign R11C32_GT00 = R20C32_GT00;
assign R11C32_GT10 = R20C32_GT10;
assign R12C32_GT00 = R20C32_GT00;
assign R12C32_GT10 = R20C32_GT10;
assign R13C32_GT00 = R20C32_GT00;
assign R13C32_GT10 = R20C32_GT10;
assign R14C32_GT00 = R20C32_GT00;
assign R14C32_GT10 = R20C32_GT10;
assign R15C32_GT00 = R20C32_GT00;
assign R15C32_GT10 = R20C32_GT10;
assign R16C32_GT00 = R20C32_GT00;
assign R16C32_GT10 = R20C32_GT10;
assign R17C32_GT00 = R20C32_GT00;
assign R17C32_GT10 = R20C32_GT10;
assign R18C32_GT00 = R20C32_GT00;
assign R18C32_GT10 = R20C32_GT10;
assign R21C32_GT00 = R20C32_GT00;
assign R21C32_GT10 = R20C32_GT10;
assign R22C32_GT00 = R20C32_GT00;
assign R22C32_GT10 = R20C32_GT10;
assign R23C32_GT00 = R20C32_GT00;
assign R23C32_GT10 = R20C32_GT10;
assign R24C32_GT00 = R20C32_GT00;
assign R24C32_GT10 = R20C32_GT10;
assign R25C32_GT00 = R20C32_GT00;
assign R25C32_GT10 = R20C32_GT10;
assign R26C32_GT00 = R20C32_GT00;
assign R26C32_GT10 = R20C32_GT10;
assign R27C32_GT00 = R20C32_GT00;
assign R27C32_GT10 = R20C32_GT10;
assign R2C2_GB00 = R2C4_GBO0;
assign R2C3_GB00 = R2C4_GBO0;
assign R2C4_GB00 = R2C4_GBO0;
assign R2C5_GB00 = R2C4_GBO0;
assign R2C6_GB00 = R2C4_GBO0;
assign R3C2_GB00 = R3C4_GBO0;
assign R3C3_GB00 = R3C4_GBO0;
assign R3C4_GB00 = R3C4_GBO0;
assign R3C5_GB00 = R3C4_GBO0;
assign R3C6_GB00 = R3C4_GBO0;
assign R4C2_GB00 = R4C4_GBO0;
assign R4C3_GB00 = R4C4_GBO0;
assign R4C4_GB00 = R4C4_GBO0;
assign R4C5_GB00 = R4C4_GBO0;
assign R4C6_GB00 = R4C4_GBO0;
assign R5C2_GB00 = R5C4_GBO0;
assign R5C3_GB00 = R5C4_GBO0;
assign R5C4_GB00 = R5C4_GBO0;
assign R5C5_GB00 = R5C4_GBO0;
assign R5C6_GB00 = R5C4_GBO0;
assign R6C2_GB00 = R6C4_GBO0;
assign R6C3_GB00 = R6C4_GBO0;
assign R6C4_GB00 = R6C4_GBO0;
assign R6C5_GB00 = R6C4_GBO0;
assign R6C6_GB00 = R6C4_GBO0;
assign R7C2_GB00 = R7C4_GBO0;
assign R7C3_GB00 = R7C4_GBO0;
assign R7C4_GB00 = R7C4_GBO0;
assign R7C5_GB00 = R7C4_GBO0;
assign R7C6_GB00 = R7C4_GBO0;
assign R8C2_GB00 = R8C4_GBO0;
assign R8C3_GB00 = R8C4_GBO0;
assign R8C4_GB00 = R8C4_GBO0;
assign R8C5_GB00 = R8C4_GBO0;
assign R8C6_GB00 = R8C4_GBO0;
assign R9C2_GB00 = R9C4_GBO0;
assign R9C3_GB00 = R9C4_GBO0;
assign R9C4_GB00 = R9C4_GBO0;
assign R9C5_GB00 = R9C4_GBO0;
assign R9C6_GB00 = R9C4_GBO0;
assign R2C9_GB00 = R2C8_GBO0;
assign R2C10_GB00 = R2C8_GBO0;
assign R2C7_GB00 = R2C8_GBO0;
assign R2C8_GB00 = R2C8_GBO0;
assign R3C9_GB00 = R3C8_GBO0;
assign R3C10_GB00 = R3C8_GBO0;
assign R3C7_GB00 = R3C8_GBO0;
assign R3C8_GB00 = R3C8_GBO0;
assign R4C9_GB00 = R4C8_GBO0;
assign R4C10_GB00 = R4C8_GBO0;
assign R4C7_GB00 = R4C8_GBO0;
assign R4C8_GB00 = R4C8_GBO0;
assign R5C9_GB00 = R5C8_GBO0;
assign R5C10_GB00 = R5C8_GBO0;
assign R5C7_GB00 = R5C8_GBO0;
assign R5C8_GB00 = R5C8_GBO0;
assign R6C9_GB00 = R6C8_GBO0;
assign R6C10_GB00 = R6C8_GBO0;
assign R6C7_GB00 = R6C8_GBO0;
assign R6C8_GB00 = R6C8_GBO0;
assign R7C9_GB00 = R7C8_GBO0;
assign R7C10_GB00 = R7C8_GBO0;
assign R7C7_GB00 = R7C8_GBO0;
assign R7C8_GB00 = R7C8_GBO0;
assign R8C9_GB00 = R8C8_GBO0;
assign R8C10_GB00 = R8C8_GBO0;
assign R8C7_GB00 = R8C8_GBO0;
assign R8C8_GB00 = R8C8_GBO0;
assign R9C9_GB00 = R9C8_GBO0;
assign R9C10_GB00 = R9C8_GBO0;
assign R9C7_GB00 = R9C8_GBO0;
assign R9C8_GB00 = R9C8_GBO0;
assign R2C11_GB00 = R2C12_GBO0;
assign R2C12_GB00 = R2C12_GBO0;
assign R2C13_GB00 = R2C12_GBO0;
assign R2C14_GB00 = R2C12_GBO0;
assign R3C11_GB00 = R3C12_GBO0;
assign R3C12_GB00 = R3C12_GBO0;
assign R3C13_GB00 = R3C12_GBO0;
assign R3C14_GB00 = R3C12_GBO0;
assign R4C11_GB00 = R4C12_GBO0;
assign R4C12_GB00 = R4C12_GBO0;
assign R4C13_GB00 = R4C12_GBO0;
assign R4C14_GB00 = R4C12_GBO0;
assign R5C11_GB00 = R5C12_GBO0;
assign R5C12_GB00 = R5C12_GBO0;
assign R5C13_GB00 = R5C12_GBO0;
assign R5C14_GB00 = R5C12_GBO0;
assign R6C11_GB00 = R6C12_GBO0;
assign R6C12_GB00 = R6C12_GBO0;
assign R6C13_GB00 = R6C12_GBO0;
assign R6C14_GB00 = R6C12_GBO0;
assign R7C11_GB00 = R7C12_GBO0;
assign R7C12_GB00 = R7C12_GBO0;
assign R7C13_GB00 = R7C12_GBO0;
assign R7C14_GB00 = R7C12_GBO0;
assign R8C11_GB00 = R8C12_GBO0;
assign R8C12_GB00 = R8C12_GBO0;
assign R8C13_GB00 = R8C12_GBO0;
assign R8C14_GB00 = R8C12_GBO0;
assign R9C11_GB00 = R9C12_GBO0;
assign R9C12_GB00 = R9C12_GBO0;
assign R9C13_GB00 = R9C12_GBO0;
assign R9C14_GB00 = R9C12_GBO0;
assign R2C17_GB00 = R2C16_GBO0;
assign R2C18_GB00 = R2C16_GBO0;
assign R2C15_GB00 = R2C16_GBO0;
assign R2C16_GB00 = R2C16_GBO0;
assign R3C17_GB00 = R3C16_GBO0;
assign R3C18_GB00 = R3C16_GBO0;
assign R3C15_GB00 = R3C16_GBO0;
assign R3C16_GB00 = R3C16_GBO0;
assign R4C17_GB00 = R4C16_GBO0;
assign R4C18_GB00 = R4C16_GBO0;
assign R4C15_GB00 = R4C16_GBO0;
assign R4C16_GB00 = R4C16_GBO0;
assign R5C17_GB00 = R5C16_GBO0;
assign R5C18_GB00 = R5C16_GBO0;
assign R5C15_GB00 = R5C16_GBO0;
assign R5C16_GB00 = R5C16_GBO0;
assign R6C17_GB00 = R6C16_GBO0;
assign R6C18_GB00 = R6C16_GBO0;
assign R6C15_GB00 = R6C16_GBO0;
assign R6C16_GB00 = R6C16_GBO0;
assign R7C17_GB00 = R7C16_GBO0;
assign R7C18_GB00 = R7C16_GBO0;
assign R7C15_GB00 = R7C16_GBO0;
assign R7C16_GB00 = R7C16_GBO0;
assign R8C17_GB00 = R8C16_GBO0;
assign R8C18_GB00 = R8C16_GBO0;
assign R8C15_GB00 = R8C16_GBO0;
assign R8C16_GB00 = R8C16_GBO0;
assign R9C17_GB00 = R9C16_GBO0;
assign R9C18_GB00 = R9C16_GBO0;
assign R9C15_GB00 = R9C16_GBO0;
assign R9C16_GB00 = R9C16_GBO0;
assign R2C19_GB00 = R2C20_GBO0;
assign R2C20_GB00 = R2C20_GBO0;
assign R2C21_GB00 = R2C20_GBO0;
assign R2C22_GB00 = R2C20_GBO0;
assign R3C19_GB00 = R3C20_GBO0;
assign R3C20_GB00 = R3C20_GBO0;
assign R3C21_GB00 = R3C20_GBO0;
assign R3C22_GB00 = R3C20_GBO0;
assign R4C19_GB00 = R4C20_GBO0;
assign R4C20_GB00 = R4C20_GBO0;
assign R4C21_GB00 = R4C20_GBO0;
assign R4C22_GB00 = R4C20_GBO0;
assign R5C19_GB00 = R5C20_GBO0;
assign R5C20_GB00 = R5C20_GBO0;
assign R5C21_GB00 = R5C20_GBO0;
assign R5C22_GB00 = R5C20_GBO0;
assign R6C19_GB00 = R6C20_GBO0;
assign R6C20_GB00 = R6C20_GBO0;
assign R6C21_GB00 = R6C20_GBO0;
assign R6C22_GB00 = R6C20_GBO0;
assign R7C19_GB00 = R7C20_GBO0;
assign R7C20_GB00 = R7C20_GBO0;
assign R7C21_GB00 = R7C20_GBO0;
assign R7C22_GB00 = R7C20_GBO0;
assign R8C19_GB00 = R8C20_GBO0;
assign R8C20_GB00 = R8C20_GBO0;
assign R8C21_GB00 = R8C20_GBO0;
assign R8C22_GB00 = R8C20_GBO0;
assign R9C19_GB00 = R9C20_GBO0;
assign R9C20_GB00 = R9C20_GBO0;
assign R9C21_GB00 = R9C20_GBO0;
assign R9C22_GB00 = R9C20_GBO0;
assign R2C23_GB00 = R2C24_GBO0;
assign R2C24_GB00 = R2C24_GBO0;
assign R2C25_GB00 = R2C24_GBO0;
assign R2C26_GB00 = R2C24_GBO0;
assign R2C27_GB00 = R2C24_GBO0;
assign R2C28_GB00 = R2C24_GBO0;
assign R3C23_GB00 = R3C24_GBO0;
assign R3C24_GB00 = R3C24_GBO0;
assign R3C25_GB00 = R3C24_GBO0;
assign R3C26_GB00 = R3C24_GBO0;
assign R3C27_GB00 = R3C24_GBO0;
assign R3C28_GB00 = R3C24_GBO0;
assign R4C23_GB00 = R4C24_GBO0;
assign R4C24_GB00 = R4C24_GBO0;
assign R4C25_GB00 = R4C24_GBO0;
assign R4C26_GB00 = R4C24_GBO0;
assign R4C27_GB00 = R4C24_GBO0;
assign R4C28_GB00 = R4C24_GBO0;
assign R5C23_GB00 = R5C24_GBO0;
assign R5C24_GB00 = R5C24_GBO0;
assign R5C25_GB00 = R5C24_GBO0;
assign R5C26_GB00 = R5C24_GBO0;
assign R5C27_GB00 = R5C24_GBO0;
assign R5C28_GB00 = R5C24_GBO0;
assign R6C23_GB00 = R6C24_GBO0;
assign R6C24_GB00 = R6C24_GBO0;
assign R6C25_GB00 = R6C24_GBO0;
assign R6C26_GB00 = R6C24_GBO0;
assign R6C27_GB00 = R6C24_GBO0;
assign R6C28_GB00 = R6C24_GBO0;
assign R7C23_GB00 = R7C24_GBO0;
assign R7C24_GB00 = R7C24_GBO0;
assign R7C25_GB00 = R7C24_GBO0;
assign R7C26_GB00 = R7C24_GBO0;
assign R7C27_GB00 = R7C24_GBO0;
assign R7C28_GB00 = R7C24_GBO0;
assign R8C23_GB00 = R8C24_GBO0;
assign R8C24_GB00 = R8C24_GBO0;
assign R8C25_GB00 = R8C24_GBO0;
assign R8C26_GB00 = R8C24_GBO0;
assign R8C27_GB00 = R8C24_GBO0;
assign R8C28_GB00 = R8C24_GBO0;
assign R9C23_GB00 = R9C24_GBO0;
assign R9C24_GB00 = R9C24_GBO0;
assign R9C25_GB00 = R9C24_GBO0;
assign R9C26_GB00 = R9C24_GBO0;
assign R9C27_GB00 = R9C24_GBO0;
assign R9C28_GB00 = R9C24_GBO0;
assign R2C2_GB10 = R2C3_GBO0;
assign R2C3_GB10 = R2C3_GBO0;
assign R2C4_GB10 = R2C3_GBO0;
assign R2C5_GB10 = R2C3_GBO0;
assign R3C2_GB10 = R3C3_GBO0;
assign R3C3_GB10 = R3C3_GBO0;
assign R3C4_GB10 = R3C3_GBO0;
assign R3C5_GB10 = R3C3_GBO0;
assign R4C2_GB10 = R4C3_GBO0;
assign R4C3_GB10 = R4C3_GBO0;
assign R4C4_GB10 = R4C3_GBO0;
assign R4C5_GB10 = R4C3_GBO0;
assign R5C2_GB10 = R5C3_GBO0;
assign R5C3_GB10 = R5C3_GBO0;
assign R5C4_GB10 = R5C3_GBO0;
assign R5C5_GB10 = R5C3_GBO0;
assign R6C2_GB10 = R6C3_GBO0;
assign R6C3_GB10 = R6C3_GBO0;
assign R6C4_GB10 = R6C3_GBO0;
assign R6C5_GB10 = R6C3_GBO0;
assign R7C2_GB10 = R7C3_GBO0;
assign R7C3_GB10 = R7C3_GBO0;
assign R7C4_GB10 = R7C3_GBO0;
assign R7C5_GB10 = R7C3_GBO0;
assign R8C2_GB10 = R8C3_GBO0;
assign R8C3_GB10 = R8C3_GBO0;
assign R8C4_GB10 = R8C3_GBO0;
assign R8C5_GB10 = R8C3_GBO0;
assign R9C2_GB10 = R9C3_GBO0;
assign R9C3_GB10 = R9C3_GBO0;
assign R9C4_GB10 = R9C3_GBO0;
assign R9C5_GB10 = R9C3_GBO0;
assign R2C9_GB10 = R2C7_GBO0;
assign R2C6_GB10 = R2C7_GBO0;
assign R2C7_GB10 = R2C7_GBO0;
assign R2C8_GB10 = R2C7_GBO0;
assign R3C9_GB10 = R3C7_GBO0;
assign R3C6_GB10 = R3C7_GBO0;
assign R3C7_GB10 = R3C7_GBO0;
assign R3C8_GB10 = R3C7_GBO0;
assign R4C9_GB10 = R4C7_GBO0;
assign R4C6_GB10 = R4C7_GBO0;
assign R4C7_GB10 = R4C7_GBO0;
assign R4C8_GB10 = R4C7_GBO0;
assign R5C9_GB10 = R5C7_GBO0;
assign R5C6_GB10 = R5C7_GBO0;
assign R5C7_GB10 = R5C7_GBO0;
assign R5C8_GB10 = R5C7_GBO0;
assign R6C9_GB10 = R6C7_GBO0;
assign R6C6_GB10 = R6C7_GBO0;
assign R6C7_GB10 = R6C7_GBO0;
assign R6C8_GB10 = R6C7_GBO0;
assign R7C9_GB10 = R7C7_GBO0;
assign R7C6_GB10 = R7C7_GBO0;
assign R7C7_GB10 = R7C7_GBO0;
assign R7C8_GB10 = R7C7_GBO0;
assign R8C9_GB10 = R8C7_GBO0;
assign R8C6_GB10 = R8C7_GBO0;
assign R8C7_GB10 = R8C7_GBO0;
assign R8C8_GB10 = R8C7_GBO0;
assign R9C9_GB10 = R9C7_GBO0;
assign R9C6_GB10 = R9C7_GBO0;
assign R9C7_GB10 = R9C7_GBO0;
assign R9C8_GB10 = R9C7_GBO0;
assign R2C10_GB10 = R2C11_GBO0;
assign R2C11_GB10 = R2C11_GBO0;
assign R2C12_GB10 = R2C11_GBO0;
assign R2C13_GB10 = R2C11_GBO0;
assign R3C10_GB10 = R3C11_GBO0;
assign R3C11_GB10 = R3C11_GBO0;
assign R3C12_GB10 = R3C11_GBO0;
assign R3C13_GB10 = R3C11_GBO0;
assign R4C10_GB10 = R4C11_GBO0;
assign R4C11_GB10 = R4C11_GBO0;
assign R4C12_GB10 = R4C11_GBO0;
assign R4C13_GB10 = R4C11_GBO0;
assign R5C10_GB10 = R5C11_GBO0;
assign R5C11_GB10 = R5C11_GBO0;
assign R5C12_GB10 = R5C11_GBO0;
assign R5C13_GB10 = R5C11_GBO0;
assign R6C10_GB10 = R6C11_GBO0;
assign R6C11_GB10 = R6C11_GBO0;
assign R6C12_GB10 = R6C11_GBO0;
assign R6C13_GB10 = R6C11_GBO0;
assign R7C10_GB10 = R7C11_GBO0;
assign R7C11_GB10 = R7C11_GBO0;
assign R7C12_GB10 = R7C11_GBO0;
assign R7C13_GB10 = R7C11_GBO0;
assign R8C10_GB10 = R8C11_GBO0;
assign R8C11_GB10 = R8C11_GBO0;
assign R8C12_GB10 = R8C11_GBO0;
assign R8C13_GB10 = R8C11_GBO0;
assign R9C10_GB10 = R9C11_GBO0;
assign R9C11_GB10 = R9C11_GBO0;
assign R9C12_GB10 = R9C11_GBO0;
assign R9C13_GB10 = R9C11_GBO0;
assign R2C17_GB10 = R2C15_GBO0;
assign R2C14_GB10 = R2C15_GBO0;
assign R2C15_GB10 = R2C15_GBO0;
assign R2C16_GB10 = R2C15_GBO0;
assign R3C17_GB10 = R3C15_GBO0;
assign R3C14_GB10 = R3C15_GBO0;
assign R3C15_GB10 = R3C15_GBO0;
assign R3C16_GB10 = R3C15_GBO0;
assign R4C17_GB10 = R4C15_GBO0;
assign R4C14_GB10 = R4C15_GBO0;
assign R4C15_GB10 = R4C15_GBO0;
assign R4C16_GB10 = R4C15_GBO0;
assign R5C17_GB10 = R5C15_GBO0;
assign R5C14_GB10 = R5C15_GBO0;
assign R5C15_GB10 = R5C15_GBO0;
assign R5C16_GB10 = R5C15_GBO0;
assign R6C17_GB10 = R6C15_GBO0;
assign R6C14_GB10 = R6C15_GBO0;
assign R6C15_GB10 = R6C15_GBO0;
assign R6C16_GB10 = R6C15_GBO0;
assign R7C17_GB10 = R7C15_GBO0;
assign R7C14_GB10 = R7C15_GBO0;
assign R7C15_GB10 = R7C15_GBO0;
assign R7C16_GB10 = R7C15_GBO0;
assign R8C17_GB10 = R8C15_GBO0;
assign R8C14_GB10 = R8C15_GBO0;
assign R8C15_GB10 = R8C15_GBO0;
assign R8C16_GB10 = R8C15_GBO0;
assign R9C17_GB10 = R9C15_GBO0;
assign R9C14_GB10 = R9C15_GBO0;
assign R9C15_GB10 = R9C15_GBO0;
assign R9C16_GB10 = R9C15_GBO0;
assign R2C18_GB10 = R2C19_GBO0;
assign R2C19_GB10 = R2C19_GBO0;
assign R2C20_GB10 = R2C19_GBO0;
assign R2C21_GB10 = R2C19_GBO0;
assign R3C18_GB10 = R3C19_GBO0;
assign R3C19_GB10 = R3C19_GBO0;
assign R3C20_GB10 = R3C19_GBO0;
assign R3C21_GB10 = R3C19_GBO0;
assign R4C18_GB10 = R4C19_GBO0;
assign R4C19_GB10 = R4C19_GBO0;
assign R4C20_GB10 = R4C19_GBO0;
assign R4C21_GB10 = R4C19_GBO0;
assign R5C18_GB10 = R5C19_GBO0;
assign R5C19_GB10 = R5C19_GBO0;
assign R5C20_GB10 = R5C19_GBO0;
assign R5C21_GB10 = R5C19_GBO0;
assign R6C18_GB10 = R6C19_GBO0;
assign R6C19_GB10 = R6C19_GBO0;
assign R6C20_GB10 = R6C19_GBO0;
assign R6C21_GB10 = R6C19_GBO0;
assign R7C18_GB10 = R7C19_GBO0;
assign R7C19_GB10 = R7C19_GBO0;
assign R7C20_GB10 = R7C19_GBO0;
assign R7C21_GB10 = R7C19_GBO0;
assign R8C18_GB10 = R8C19_GBO0;
assign R8C19_GB10 = R8C19_GBO0;
assign R8C20_GB10 = R8C19_GBO0;
assign R8C21_GB10 = R8C19_GBO0;
assign R9C18_GB10 = R9C19_GBO0;
assign R9C19_GB10 = R9C19_GBO0;
assign R9C20_GB10 = R9C19_GBO0;
assign R9C21_GB10 = R9C19_GBO0;
assign R2C25_GB10 = R2C23_GBO0;
assign R2C22_GB10 = R2C23_GBO0;
assign R2C23_GB10 = R2C23_GBO0;
assign R2C24_GB10 = R2C23_GBO0;
assign R3C25_GB10 = R3C23_GBO0;
assign R3C22_GB10 = R3C23_GBO0;
assign R3C23_GB10 = R3C23_GBO0;
assign R3C24_GB10 = R3C23_GBO0;
assign R4C25_GB10 = R4C23_GBO0;
assign R4C22_GB10 = R4C23_GBO0;
assign R4C23_GB10 = R4C23_GBO0;
assign R4C24_GB10 = R4C23_GBO0;
assign R5C25_GB10 = R5C23_GBO0;
assign R5C22_GB10 = R5C23_GBO0;
assign R5C23_GB10 = R5C23_GBO0;
assign R5C24_GB10 = R5C23_GBO0;
assign R6C25_GB10 = R6C23_GBO0;
assign R6C22_GB10 = R6C23_GBO0;
assign R6C23_GB10 = R6C23_GBO0;
assign R6C24_GB10 = R6C23_GBO0;
assign R7C25_GB10 = R7C23_GBO0;
assign R7C22_GB10 = R7C23_GBO0;
assign R7C23_GB10 = R7C23_GBO0;
assign R7C24_GB10 = R7C23_GBO0;
assign R8C25_GB10 = R8C23_GBO0;
assign R8C22_GB10 = R8C23_GBO0;
assign R8C23_GB10 = R8C23_GBO0;
assign R8C24_GB10 = R8C23_GBO0;
assign R9C25_GB10 = R9C23_GBO0;
assign R9C22_GB10 = R9C23_GBO0;
assign R9C23_GB10 = R9C23_GBO0;
assign R9C24_GB10 = R9C23_GBO0;
assign R2C26_GB10 = R2C27_GBO0;
assign R2C27_GB10 = R2C27_GBO0;
assign R2C28_GB10 = R2C27_GBO0;
assign R3C26_GB10 = R3C27_GBO0;
assign R3C27_GB10 = R3C27_GBO0;
assign R3C28_GB10 = R3C27_GBO0;
assign R4C26_GB10 = R4C27_GBO0;
assign R4C27_GB10 = R4C27_GBO0;
assign R4C28_GB10 = R4C27_GBO0;
assign R5C26_GB10 = R5C27_GBO0;
assign R5C27_GB10 = R5C27_GBO0;
assign R5C28_GB10 = R5C27_GBO0;
assign R6C26_GB10 = R6C27_GBO0;
assign R6C27_GB10 = R6C27_GBO0;
assign R6C28_GB10 = R6C27_GBO0;
assign R7C26_GB10 = R7C27_GBO0;
assign R7C27_GB10 = R7C27_GBO0;
assign R7C28_GB10 = R7C27_GBO0;
assign R8C26_GB10 = R8C27_GBO0;
assign R8C27_GB10 = R8C27_GBO0;
assign R8C28_GB10 = R8C27_GBO0;
assign R9C26_GB10 = R9C27_GBO0;
assign R9C27_GB10 = R9C27_GBO0;
assign R9C28_GB10 = R9C27_GBO0;
assign R2C2_GB20 = R2C2_GBO0;
assign R2C3_GB20 = R2C2_GBO0;
assign R2C4_GB20 = R2C2_GBO0;
assign R3C2_GB20 = R3C2_GBO0;
assign R3C3_GB20 = R3C2_GBO0;
assign R3C4_GB20 = R3C2_GBO0;
assign R4C2_GB20 = R4C2_GBO0;
assign R4C3_GB20 = R4C2_GBO0;
assign R4C4_GB20 = R4C2_GBO0;
assign R5C2_GB20 = R5C2_GBO0;
assign R5C3_GB20 = R5C2_GBO0;
assign R5C4_GB20 = R5C2_GBO0;
assign R6C2_GB20 = R6C2_GBO0;
assign R6C3_GB20 = R6C2_GBO0;
assign R6C4_GB20 = R6C2_GBO0;
assign R7C2_GB20 = R7C2_GBO0;
assign R7C3_GB20 = R7C2_GBO0;
assign R7C4_GB20 = R7C2_GBO0;
assign R8C2_GB20 = R8C2_GBO0;
assign R8C3_GB20 = R8C2_GBO0;
assign R8C4_GB20 = R8C2_GBO0;
assign R9C2_GB20 = R9C2_GBO0;
assign R9C3_GB20 = R9C2_GBO0;
assign R9C4_GB20 = R9C2_GBO0;
assign R2C5_GB20 = R2C6_GBO0;
assign R2C6_GB20 = R2C6_GBO0;
assign R2C7_GB20 = R2C6_GBO0;
assign R2C8_GB20 = R2C6_GBO0;
assign R3C5_GB20 = R3C6_GBO0;
assign R3C6_GB20 = R3C6_GBO0;
assign R3C7_GB20 = R3C6_GBO0;
assign R3C8_GB20 = R3C6_GBO0;
assign R4C5_GB20 = R4C6_GBO0;
assign R4C6_GB20 = R4C6_GBO0;
assign R4C7_GB20 = R4C6_GBO0;
assign R4C8_GB20 = R4C6_GBO0;
assign R5C5_GB20 = R5C6_GBO0;
assign R5C6_GB20 = R5C6_GBO0;
assign R5C7_GB20 = R5C6_GBO0;
assign R5C8_GB20 = R5C6_GBO0;
assign R6C5_GB20 = R6C6_GBO0;
assign R6C6_GB20 = R6C6_GBO0;
assign R6C7_GB20 = R6C6_GBO0;
assign R6C8_GB20 = R6C6_GBO0;
assign R7C5_GB20 = R7C6_GBO0;
assign R7C6_GB20 = R7C6_GBO0;
assign R7C7_GB20 = R7C6_GBO0;
assign R7C8_GB20 = R7C6_GBO0;
assign R8C5_GB20 = R8C6_GBO0;
assign R8C6_GB20 = R8C6_GBO0;
assign R8C7_GB20 = R8C6_GBO0;
assign R8C8_GB20 = R8C6_GBO0;
assign R9C5_GB20 = R9C6_GBO0;
assign R9C6_GB20 = R9C6_GBO0;
assign R9C7_GB20 = R9C6_GBO0;
assign R9C8_GB20 = R9C6_GBO0;
assign R2C9_GB20 = R2C10_GBO0;
assign R2C10_GB20 = R2C10_GBO0;
assign R2C11_GB20 = R2C10_GBO0;
assign R2C12_GB20 = R2C10_GBO0;
assign R3C9_GB20 = R3C10_GBO0;
assign R3C10_GB20 = R3C10_GBO0;
assign R3C11_GB20 = R3C10_GBO0;
assign R3C12_GB20 = R3C10_GBO0;
assign R4C9_GB20 = R4C10_GBO0;
assign R4C10_GB20 = R4C10_GBO0;
assign R4C11_GB20 = R4C10_GBO0;
assign R4C12_GB20 = R4C10_GBO0;
assign R5C9_GB20 = R5C10_GBO0;
assign R5C10_GB20 = R5C10_GBO0;
assign R5C11_GB20 = R5C10_GBO0;
assign R5C12_GB20 = R5C10_GBO0;
assign R6C9_GB20 = R6C10_GBO0;
assign R6C10_GB20 = R6C10_GBO0;
assign R6C11_GB20 = R6C10_GBO0;
assign R6C12_GB20 = R6C10_GBO0;
assign R7C9_GB20 = R7C10_GBO0;
assign R7C10_GB20 = R7C10_GBO0;
assign R7C11_GB20 = R7C10_GBO0;
assign R7C12_GB20 = R7C10_GBO0;
assign R8C9_GB20 = R8C10_GBO0;
assign R8C10_GB20 = R8C10_GBO0;
assign R8C11_GB20 = R8C10_GBO0;
assign R8C12_GB20 = R8C10_GBO0;
assign R9C9_GB20 = R9C10_GBO0;
assign R9C10_GB20 = R9C10_GBO0;
assign R9C11_GB20 = R9C10_GBO0;
assign R9C12_GB20 = R9C10_GBO0;
assign R2C13_GB20 = R2C14_GBO0;
assign R2C14_GB20 = R2C14_GBO0;
assign R2C15_GB20 = R2C14_GBO0;
assign R2C16_GB20 = R2C14_GBO0;
assign R3C13_GB20 = R3C14_GBO0;
assign R3C14_GB20 = R3C14_GBO0;
assign R3C15_GB20 = R3C14_GBO0;
assign R3C16_GB20 = R3C14_GBO0;
assign R4C13_GB20 = R4C14_GBO0;
assign R4C14_GB20 = R4C14_GBO0;
assign R4C15_GB20 = R4C14_GBO0;
assign R4C16_GB20 = R4C14_GBO0;
assign R5C13_GB20 = R5C14_GBO0;
assign R5C14_GB20 = R5C14_GBO0;
assign R5C15_GB20 = R5C14_GBO0;
assign R5C16_GB20 = R5C14_GBO0;
assign R6C13_GB20 = R6C14_GBO0;
assign R6C14_GB20 = R6C14_GBO0;
assign R6C15_GB20 = R6C14_GBO0;
assign R6C16_GB20 = R6C14_GBO0;
assign R7C13_GB20 = R7C14_GBO0;
assign R7C14_GB20 = R7C14_GBO0;
assign R7C15_GB20 = R7C14_GBO0;
assign R7C16_GB20 = R7C14_GBO0;
assign R8C13_GB20 = R8C14_GBO0;
assign R8C14_GB20 = R8C14_GBO0;
assign R8C15_GB20 = R8C14_GBO0;
assign R8C16_GB20 = R8C14_GBO0;
assign R9C13_GB20 = R9C14_GBO0;
assign R9C14_GB20 = R9C14_GBO0;
assign R9C15_GB20 = R9C14_GBO0;
assign R9C16_GB20 = R9C14_GBO0;
assign R2C17_GB20 = R2C18_GBO0;
assign R2C18_GB20 = R2C18_GBO0;
assign R2C19_GB20 = R2C18_GBO0;
assign R2C20_GB20 = R2C18_GBO0;
assign R3C17_GB20 = R3C18_GBO0;
assign R3C18_GB20 = R3C18_GBO0;
assign R3C19_GB20 = R3C18_GBO0;
assign R3C20_GB20 = R3C18_GBO0;
assign R4C17_GB20 = R4C18_GBO0;
assign R4C18_GB20 = R4C18_GBO0;
assign R4C19_GB20 = R4C18_GBO0;
assign R4C20_GB20 = R4C18_GBO0;
assign R5C17_GB20 = R5C18_GBO0;
assign R5C18_GB20 = R5C18_GBO0;
assign R5C19_GB20 = R5C18_GBO0;
assign R5C20_GB20 = R5C18_GBO0;
assign R6C17_GB20 = R6C18_GBO0;
assign R6C18_GB20 = R6C18_GBO0;
assign R6C19_GB20 = R6C18_GBO0;
assign R6C20_GB20 = R6C18_GBO0;
assign R7C17_GB20 = R7C18_GBO0;
assign R7C18_GB20 = R7C18_GBO0;
assign R7C19_GB20 = R7C18_GBO0;
assign R7C20_GB20 = R7C18_GBO0;
assign R8C17_GB20 = R8C18_GBO0;
assign R8C18_GB20 = R8C18_GBO0;
assign R8C19_GB20 = R8C18_GBO0;
assign R8C20_GB20 = R8C18_GBO0;
assign R9C17_GB20 = R9C18_GBO0;
assign R9C18_GB20 = R9C18_GBO0;
assign R9C19_GB20 = R9C18_GBO0;
assign R9C20_GB20 = R9C18_GBO0;
assign R2C21_GB20 = R2C22_GBO0;
assign R2C22_GB20 = R2C22_GBO0;
assign R2C23_GB20 = R2C22_GBO0;
assign R2C24_GB20 = R2C22_GBO0;
assign R3C21_GB20 = R3C22_GBO0;
assign R3C22_GB20 = R3C22_GBO0;
assign R3C23_GB20 = R3C22_GBO0;
assign R3C24_GB20 = R3C22_GBO0;
assign R4C21_GB20 = R4C22_GBO0;
assign R4C22_GB20 = R4C22_GBO0;
assign R4C23_GB20 = R4C22_GBO0;
assign R4C24_GB20 = R4C22_GBO0;
assign R5C21_GB20 = R5C22_GBO0;
assign R5C22_GB20 = R5C22_GBO0;
assign R5C23_GB20 = R5C22_GBO0;
assign R5C24_GB20 = R5C22_GBO0;
assign R6C21_GB20 = R6C22_GBO0;
assign R6C22_GB20 = R6C22_GBO0;
assign R6C23_GB20 = R6C22_GBO0;
assign R6C24_GB20 = R6C22_GBO0;
assign R7C21_GB20 = R7C22_GBO0;
assign R7C22_GB20 = R7C22_GBO0;
assign R7C23_GB20 = R7C22_GBO0;
assign R7C24_GB20 = R7C22_GBO0;
assign R8C21_GB20 = R8C22_GBO0;
assign R8C22_GB20 = R8C22_GBO0;
assign R8C23_GB20 = R8C22_GBO0;
assign R8C24_GB20 = R8C22_GBO0;
assign R9C21_GB20 = R9C22_GBO0;
assign R9C22_GB20 = R9C22_GBO0;
assign R9C23_GB20 = R9C22_GBO0;
assign R9C24_GB20 = R9C22_GBO0;
assign R2C25_GB20 = R2C26_GBO0;
assign R2C26_GB20 = R2C26_GBO0;
assign R2C27_GB20 = R2C26_GBO0;
assign R2C28_GB20 = R2C26_GBO0;
assign R3C25_GB20 = R3C26_GBO0;
assign R3C26_GB20 = R3C26_GBO0;
assign R3C27_GB20 = R3C26_GBO0;
assign R3C28_GB20 = R3C26_GBO0;
assign R4C25_GB20 = R4C26_GBO0;
assign R4C26_GB20 = R4C26_GBO0;
assign R4C27_GB20 = R4C26_GBO0;
assign R4C28_GB20 = R4C26_GBO0;
assign R5C25_GB20 = R5C26_GBO0;
assign R5C26_GB20 = R5C26_GBO0;
assign R5C27_GB20 = R5C26_GBO0;
assign R5C28_GB20 = R5C26_GBO0;
assign R6C25_GB20 = R6C26_GBO0;
assign R6C26_GB20 = R6C26_GBO0;
assign R6C27_GB20 = R6C26_GBO0;
assign R6C28_GB20 = R6C26_GBO0;
assign R7C25_GB20 = R7C26_GBO0;
assign R7C26_GB20 = R7C26_GBO0;
assign R7C27_GB20 = R7C26_GBO0;
assign R7C28_GB20 = R7C26_GBO0;
assign R8C25_GB20 = R8C26_GBO0;
assign R8C26_GB20 = R8C26_GBO0;
assign R8C27_GB20 = R8C26_GBO0;
assign R8C28_GB20 = R8C26_GBO0;
assign R9C25_GB20 = R9C26_GBO0;
assign R9C26_GB20 = R9C26_GBO0;
assign R9C27_GB20 = R9C26_GBO0;
assign R9C28_GB20 = R9C26_GBO0;
assign R2C2_GB30 = R2C1_GBO0;
assign R2C3_GB30 = R2C1_GBO0;
assign R3C2_GB30 = R3C1_GBO0;
assign R3C3_GB30 = R3C1_GBO0;
assign R4C2_GB30 = R4C1_GBO0;
assign R4C3_GB30 = R4C1_GBO0;
assign R5C2_GB30 = R5C1_GBO0;
assign R5C3_GB30 = R5C1_GBO0;
assign R6C2_GB30 = R6C1_GBO0;
assign R6C3_GB30 = R6C1_GBO0;
assign R7C2_GB30 = R7C1_GBO0;
assign R7C3_GB30 = R7C1_GBO0;
assign R8C2_GB30 = R8C1_GBO0;
assign R8C3_GB30 = R8C1_GBO0;
assign R9C2_GB30 = R9C1_GBO0;
assign R9C3_GB30 = R9C1_GBO0;
assign R2C4_GB30 = R2C5_GBO0;
assign R2C5_GB30 = R2C5_GBO0;
assign R2C6_GB30 = R2C5_GBO0;
assign R2C7_GB30 = R2C5_GBO0;
assign R3C4_GB30 = R3C5_GBO0;
assign R3C5_GB30 = R3C5_GBO0;
assign R3C6_GB30 = R3C5_GBO0;
assign R3C7_GB30 = R3C5_GBO0;
assign R4C4_GB30 = R4C5_GBO0;
assign R4C5_GB30 = R4C5_GBO0;
assign R4C6_GB30 = R4C5_GBO0;
assign R4C7_GB30 = R4C5_GBO0;
assign R5C4_GB30 = R5C5_GBO0;
assign R5C5_GB30 = R5C5_GBO0;
assign R5C6_GB30 = R5C5_GBO0;
assign R5C7_GB30 = R5C5_GBO0;
assign R6C4_GB30 = R6C5_GBO0;
assign R6C5_GB30 = R6C5_GBO0;
assign R6C6_GB30 = R6C5_GBO0;
assign R6C7_GB30 = R6C5_GBO0;
assign R7C4_GB30 = R7C5_GBO0;
assign R7C5_GB30 = R7C5_GBO0;
assign R7C6_GB30 = R7C5_GBO0;
assign R7C7_GB30 = R7C5_GBO0;
assign R8C4_GB30 = R8C5_GBO0;
assign R8C5_GB30 = R8C5_GBO0;
assign R8C6_GB30 = R8C5_GBO0;
assign R8C7_GB30 = R8C5_GBO0;
assign R9C4_GB30 = R9C5_GBO0;
assign R9C5_GB30 = R9C5_GBO0;
assign R9C6_GB30 = R9C5_GBO0;
assign R9C7_GB30 = R9C5_GBO0;
assign R2C9_GB30 = R2C9_GBO0;
assign R2C10_GB30 = R2C9_GBO0;
assign R2C11_GB30 = R2C9_GBO0;
assign R2C8_GB30 = R2C9_GBO0;
assign R3C9_GB30 = R3C9_GBO0;
assign R3C10_GB30 = R3C9_GBO0;
assign R3C11_GB30 = R3C9_GBO0;
assign R3C8_GB30 = R3C9_GBO0;
assign R4C9_GB30 = R4C9_GBO0;
assign R4C10_GB30 = R4C9_GBO0;
assign R4C11_GB30 = R4C9_GBO0;
assign R4C8_GB30 = R4C9_GBO0;
assign R5C9_GB30 = R5C9_GBO0;
assign R5C10_GB30 = R5C9_GBO0;
assign R5C11_GB30 = R5C9_GBO0;
assign R5C8_GB30 = R5C9_GBO0;
assign R6C9_GB30 = R6C9_GBO0;
assign R6C10_GB30 = R6C9_GBO0;
assign R6C11_GB30 = R6C9_GBO0;
assign R6C8_GB30 = R6C9_GBO0;
assign R7C9_GB30 = R7C9_GBO0;
assign R7C10_GB30 = R7C9_GBO0;
assign R7C11_GB30 = R7C9_GBO0;
assign R7C8_GB30 = R7C9_GBO0;
assign R8C9_GB30 = R8C9_GBO0;
assign R8C10_GB30 = R8C9_GBO0;
assign R8C11_GB30 = R8C9_GBO0;
assign R8C8_GB30 = R8C9_GBO0;
assign R9C9_GB30 = R9C9_GBO0;
assign R9C10_GB30 = R9C9_GBO0;
assign R9C11_GB30 = R9C9_GBO0;
assign R9C8_GB30 = R9C9_GBO0;
assign R2C12_GB30 = R2C13_GBO0;
assign R2C13_GB30 = R2C13_GBO0;
assign R2C14_GB30 = R2C13_GBO0;
assign R2C15_GB30 = R2C13_GBO0;
assign R3C12_GB30 = R3C13_GBO0;
assign R3C13_GB30 = R3C13_GBO0;
assign R3C14_GB30 = R3C13_GBO0;
assign R3C15_GB30 = R3C13_GBO0;
assign R4C12_GB30 = R4C13_GBO0;
assign R4C13_GB30 = R4C13_GBO0;
assign R4C14_GB30 = R4C13_GBO0;
assign R4C15_GB30 = R4C13_GBO0;
assign R5C12_GB30 = R5C13_GBO0;
assign R5C13_GB30 = R5C13_GBO0;
assign R5C14_GB30 = R5C13_GBO0;
assign R5C15_GB30 = R5C13_GBO0;
assign R6C12_GB30 = R6C13_GBO0;
assign R6C13_GB30 = R6C13_GBO0;
assign R6C14_GB30 = R6C13_GBO0;
assign R6C15_GB30 = R6C13_GBO0;
assign R7C12_GB30 = R7C13_GBO0;
assign R7C13_GB30 = R7C13_GBO0;
assign R7C14_GB30 = R7C13_GBO0;
assign R7C15_GB30 = R7C13_GBO0;
assign R8C12_GB30 = R8C13_GBO0;
assign R8C13_GB30 = R8C13_GBO0;
assign R8C14_GB30 = R8C13_GBO0;
assign R8C15_GB30 = R8C13_GBO0;
assign R9C12_GB30 = R9C13_GBO0;
assign R9C13_GB30 = R9C13_GBO0;
assign R9C14_GB30 = R9C13_GBO0;
assign R9C15_GB30 = R9C13_GBO0;
assign R2C17_GB30 = R2C17_GBO0;
assign R2C18_GB30 = R2C17_GBO0;
assign R2C19_GB30 = R2C17_GBO0;
assign R2C16_GB30 = R2C17_GBO0;
assign R3C17_GB30 = R3C17_GBO0;
assign R3C18_GB30 = R3C17_GBO0;
assign R3C19_GB30 = R3C17_GBO0;
assign R3C16_GB30 = R3C17_GBO0;
assign R4C17_GB30 = R4C17_GBO0;
assign R4C18_GB30 = R4C17_GBO0;
assign R4C19_GB30 = R4C17_GBO0;
assign R4C16_GB30 = R4C17_GBO0;
assign R5C17_GB30 = R5C17_GBO0;
assign R5C18_GB30 = R5C17_GBO0;
assign R5C19_GB30 = R5C17_GBO0;
assign R5C16_GB30 = R5C17_GBO0;
assign R6C17_GB30 = R6C17_GBO0;
assign R6C18_GB30 = R6C17_GBO0;
assign R6C19_GB30 = R6C17_GBO0;
assign R6C16_GB30 = R6C17_GBO0;
assign R7C17_GB30 = R7C17_GBO0;
assign R7C18_GB30 = R7C17_GBO0;
assign R7C19_GB30 = R7C17_GBO0;
assign R7C16_GB30 = R7C17_GBO0;
assign R8C17_GB30 = R8C17_GBO0;
assign R8C18_GB30 = R8C17_GBO0;
assign R8C19_GB30 = R8C17_GBO0;
assign R8C16_GB30 = R8C17_GBO0;
assign R9C17_GB30 = R9C17_GBO0;
assign R9C18_GB30 = R9C17_GBO0;
assign R9C19_GB30 = R9C17_GBO0;
assign R9C16_GB30 = R9C17_GBO0;
assign R2C20_GB30 = R2C21_GBO0;
assign R2C21_GB30 = R2C21_GBO0;
assign R2C22_GB30 = R2C21_GBO0;
assign R2C23_GB30 = R2C21_GBO0;
assign R3C20_GB30 = R3C21_GBO0;
assign R3C21_GB30 = R3C21_GBO0;
assign R3C22_GB30 = R3C21_GBO0;
assign R3C23_GB30 = R3C21_GBO0;
assign R4C20_GB30 = R4C21_GBO0;
assign R4C21_GB30 = R4C21_GBO0;
assign R4C22_GB30 = R4C21_GBO0;
assign R4C23_GB30 = R4C21_GBO0;
assign R5C20_GB30 = R5C21_GBO0;
assign R5C21_GB30 = R5C21_GBO0;
assign R5C22_GB30 = R5C21_GBO0;
assign R5C23_GB30 = R5C21_GBO0;
assign R6C20_GB30 = R6C21_GBO0;
assign R6C21_GB30 = R6C21_GBO0;
assign R6C22_GB30 = R6C21_GBO0;
assign R6C23_GB30 = R6C21_GBO0;
assign R7C20_GB30 = R7C21_GBO0;
assign R7C21_GB30 = R7C21_GBO0;
assign R7C22_GB30 = R7C21_GBO0;
assign R7C23_GB30 = R7C21_GBO0;
assign R8C20_GB30 = R8C21_GBO0;
assign R8C21_GB30 = R8C21_GBO0;
assign R8C22_GB30 = R8C21_GBO0;
assign R8C23_GB30 = R8C21_GBO0;
assign R9C20_GB30 = R9C21_GBO0;
assign R9C21_GB30 = R9C21_GBO0;
assign R9C22_GB30 = R9C21_GBO0;
assign R9C23_GB30 = R9C21_GBO0;
assign R2C24_GB30 = R2C25_GBO0;
assign R2C25_GB30 = R2C25_GBO0;
assign R2C26_GB30 = R2C25_GBO0;
assign R2C27_GB30 = R2C25_GBO0;
assign R2C28_GB30 = R2C25_GBO0;
assign R3C24_GB30 = R3C25_GBO0;
assign R3C25_GB30 = R3C25_GBO0;
assign R3C26_GB30 = R3C25_GBO0;
assign R3C27_GB30 = R3C25_GBO0;
assign R3C28_GB30 = R3C25_GBO0;
assign R4C24_GB30 = R4C25_GBO0;
assign R4C25_GB30 = R4C25_GBO0;
assign R4C26_GB30 = R4C25_GBO0;
assign R4C27_GB30 = R4C25_GBO0;
assign R4C28_GB30 = R4C25_GBO0;
assign R5C24_GB30 = R5C25_GBO0;
assign R5C25_GB30 = R5C25_GBO0;
assign R5C26_GB30 = R5C25_GBO0;
assign R5C27_GB30 = R5C25_GBO0;
assign R5C28_GB30 = R5C25_GBO0;
assign R6C24_GB30 = R6C25_GBO0;
assign R6C25_GB30 = R6C25_GBO0;
assign R6C26_GB30 = R6C25_GBO0;
assign R6C27_GB30 = R6C25_GBO0;
assign R6C28_GB30 = R6C25_GBO0;
assign R7C24_GB30 = R7C25_GBO0;
assign R7C25_GB30 = R7C25_GBO0;
assign R7C26_GB30 = R7C25_GBO0;
assign R7C27_GB30 = R7C25_GBO0;
assign R7C28_GB30 = R7C25_GBO0;
assign R8C24_GB30 = R8C25_GBO0;
assign R8C25_GB30 = R8C25_GBO0;
assign R8C26_GB30 = R8C25_GBO0;
assign R8C27_GB30 = R8C25_GBO0;
assign R8C28_GB30 = R8C25_GBO0;
assign R9C24_GB30 = R9C25_GBO0;
assign R9C25_GB30 = R9C25_GBO0;
assign R9C26_GB30 = R9C25_GBO0;
assign R9C27_GB30 = R9C25_GBO0;
assign R9C28_GB30 = R9C25_GBO0;
assign R2C2_GB40 = R2C4_GBO1;
assign R2C3_GB40 = R2C4_GBO1;
assign R2C4_GB40 = R2C4_GBO1;
assign R2C5_GB40 = R2C4_GBO1;
assign R2C6_GB40 = R2C4_GBO1;
assign R3C2_GB40 = R3C4_GBO1;
assign R3C3_GB40 = R3C4_GBO1;
assign R3C4_GB40 = R3C4_GBO1;
assign R3C5_GB40 = R3C4_GBO1;
assign R3C6_GB40 = R3C4_GBO1;
assign R4C2_GB40 = R4C4_GBO1;
assign R4C3_GB40 = R4C4_GBO1;
assign R4C4_GB40 = R4C4_GBO1;
assign R4C5_GB40 = R4C4_GBO1;
assign R4C6_GB40 = R4C4_GBO1;
assign R5C2_GB40 = R5C4_GBO1;
assign R5C3_GB40 = R5C4_GBO1;
assign R5C4_GB40 = R5C4_GBO1;
assign R5C5_GB40 = R5C4_GBO1;
assign R5C6_GB40 = R5C4_GBO1;
assign R6C2_GB40 = R6C4_GBO1;
assign R6C3_GB40 = R6C4_GBO1;
assign R6C4_GB40 = R6C4_GBO1;
assign R6C5_GB40 = R6C4_GBO1;
assign R6C6_GB40 = R6C4_GBO1;
assign R7C2_GB40 = R7C4_GBO1;
assign R7C3_GB40 = R7C4_GBO1;
assign R7C4_GB40 = R7C4_GBO1;
assign R7C5_GB40 = R7C4_GBO1;
assign R7C6_GB40 = R7C4_GBO1;
assign R8C2_GB40 = R8C4_GBO1;
assign R8C3_GB40 = R8C4_GBO1;
assign R8C4_GB40 = R8C4_GBO1;
assign R8C5_GB40 = R8C4_GBO1;
assign R8C6_GB40 = R8C4_GBO1;
assign R9C2_GB40 = R9C4_GBO1;
assign R9C3_GB40 = R9C4_GBO1;
assign R9C4_GB40 = R9C4_GBO1;
assign R9C5_GB40 = R9C4_GBO1;
assign R9C6_GB40 = R9C4_GBO1;
assign R2C9_GB40 = R2C8_GBO1;
assign R2C10_GB40 = R2C8_GBO1;
assign R2C7_GB40 = R2C8_GBO1;
assign R2C8_GB40 = R2C8_GBO1;
assign R3C9_GB40 = R3C8_GBO1;
assign R3C10_GB40 = R3C8_GBO1;
assign R3C7_GB40 = R3C8_GBO1;
assign R3C8_GB40 = R3C8_GBO1;
assign R4C9_GB40 = R4C8_GBO1;
assign R4C10_GB40 = R4C8_GBO1;
assign R4C7_GB40 = R4C8_GBO1;
assign R4C8_GB40 = R4C8_GBO1;
assign R5C9_GB40 = R5C8_GBO1;
assign R5C10_GB40 = R5C8_GBO1;
assign R5C7_GB40 = R5C8_GBO1;
assign R5C8_GB40 = R5C8_GBO1;
assign R6C9_GB40 = R6C8_GBO1;
assign R6C10_GB40 = R6C8_GBO1;
assign R6C7_GB40 = R6C8_GBO1;
assign R6C8_GB40 = R6C8_GBO1;
assign R7C9_GB40 = R7C8_GBO1;
assign R7C10_GB40 = R7C8_GBO1;
assign R7C7_GB40 = R7C8_GBO1;
assign R7C8_GB40 = R7C8_GBO1;
assign R8C9_GB40 = R8C8_GBO1;
assign R8C10_GB40 = R8C8_GBO1;
assign R8C7_GB40 = R8C8_GBO1;
assign R8C8_GB40 = R8C8_GBO1;
assign R9C9_GB40 = R9C8_GBO1;
assign R9C10_GB40 = R9C8_GBO1;
assign R9C7_GB40 = R9C8_GBO1;
assign R9C8_GB40 = R9C8_GBO1;
assign R2C11_GB40 = R2C12_GBO1;
assign R2C12_GB40 = R2C12_GBO1;
assign R2C13_GB40 = R2C12_GBO1;
assign R2C14_GB40 = R2C12_GBO1;
assign R3C11_GB40 = R3C12_GBO1;
assign R3C12_GB40 = R3C12_GBO1;
assign R3C13_GB40 = R3C12_GBO1;
assign R3C14_GB40 = R3C12_GBO1;
assign R4C11_GB40 = R4C12_GBO1;
assign R4C12_GB40 = R4C12_GBO1;
assign R4C13_GB40 = R4C12_GBO1;
assign R4C14_GB40 = R4C12_GBO1;
assign R5C11_GB40 = R5C12_GBO1;
assign R5C12_GB40 = R5C12_GBO1;
assign R5C13_GB40 = R5C12_GBO1;
assign R5C14_GB40 = R5C12_GBO1;
assign R6C11_GB40 = R6C12_GBO1;
assign R6C12_GB40 = R6C12_GBO1;
assign R6C13_GB40 = R6C12_GBO1;
assign R6C14_GB40 = R6C12_GBO1;
assign R7C11_GB40 = R7C12_GBO1;
assign R7C12_GB40 = R7C12_GBO1;
assign R7C13_GB40 = R7C12_GBO1;
assign R7C14_GB40 = R7C12_GBO1;
assign R8C11_GB40 = R8C12_GBO1;
assign R8C12_GB40 = R8C12_GBO1;
assign R8C13_GB40 = R8C12_GBO1;
assign R8C14_GB40 = R8C12_GBO1;
assign R9C11_GB40 = R9C12_GBO1;
assign R9C12_GB40 = R9C12_GBO1;
assign R9C13_GB40 = R9C12_GBO1;
assign R9C14_GB40 = R9C12_GBO1;
assign R2C17_GB40 = R2C16_GBO1;
assign R2C18_GB40 = R2C16_GBO1;
assign R2C15_GB40 = R2C16_GBO1;
assign R2C16_GB40 = R2C16_GBO1;
assign R3C17_GB40 = R3C16_GBO1;
assign R3C18_GB40 = R3C16_GBO1;
assign R3C15_GB40 = R3C16_GBO1;
assign R3C16_GB40 = R3C16_GBO1;
assign R4C17_GB40 = R4C16_GBO1;
assign R4C18_GB40 = R4C16_GBO1;
assign R4C15_GB40 = R4C16_GBO1;
assign R4C16_GB40 = R4C16_GBO1;
assign R5C17_GB40 = R5C16_GBO1;
assign R5C18_GB40 = R5C16_GBO1;
assign R5C15_GB40 = R5C16_GBO1;
assign R5C16_GB40 = R5C16_GBO1;
assign R6C17_GB40 = R6C16_GBO1;
assign R6C18_GB40 = R6C16_GBO1;
assign R6C15_GB40 = R6C16_GBO1;
assign R6C16_GB40 = R6C16_GBO1;
assign R7C17_GB40 = R7C16_GBO1;
assign R7C18_GB40 = R7C16_GBO1;
assign R7C15_GB40 = R7C16_GBO1;
assign R7C16_GB40 = R7C16_GBO1;
assign R8C17_GB40 = R8C16_GBO1;
assign R8C18_GB40 = R8C16_GBO1;
assign R8C15_GB40 = R8C16_GBO1;
assign R8C16_GB40 = R8C16_GBO1;
assign R9C17_GB40 = R9C16_GBO1;
assign R9C18_GB40 = R9C16_GBO1;
assign R9C15_GB40 = R9C16_GBO1;
assign R9C16_GB40 = R9C16_GBO1;
assign R2C19_GB40 = R2C20_GBO1;
assign R2C20_GB40 = R2C20_GBO1;
assign R2C21_GB40 = R2C20_GBO1;
assign R2C22_GB40 = R2C20_GBO1;
assign R3C19_GB40 = R3C20_GBO1;
assign R3C20_GB40 = R3C20_GBO1;
assign R3C21_GB40 = R3C20_GBO1;
assign R3C22_GB40 = R3C20_GBO1;
assign R4C19_GB40 = R4C20_GBO1;
assign R4C20_GB40 = R4C20_GBO1;
assign R4C21_GB40 = R4C20_GBO1;
assign R4C22_GB40 = R4C20_GBO1;
assign R5C19_GB40 = R5C20_GBO1;
assign R5C20_GB40 = R5C20_GBO1;
assign R5C21_GB40 = R5C20_GBO1;
assign R5C22_GB40 = R5C20_GBO1;
assign R6C19_GB40 = R6C20_GBO1;
assign R6C20_GB40 = R6C20_GBO1;
assign R6C21_GB40 = R6C20_GBO1;
assign R6C22_GB40 = R6C20_GBO1;
assign R7C19_GB40 = R7C20_GBO1;
assign R7C20_GB40 = R7C20_GBO1;
assign R7C21_GB40 = R7C20_GBO1;
assign R7C22_GB40 = R7C20_GBO1;
assign R8C19_GB40 = R8C20_GBO1;
assign R8C20_GB40 = R8C20_GBO1;
assign R8C21_GB40 = R8C20_GBO1;
assign R8C22_GB40 = R8C20_GBO1;
assign R9C19_GB40 = R9C20_GBO1;
assign R9C20_GB40 = R9C20_GBO1;
assign R9C21_GB40 = R9C20_GBO1;
assign R9C22_GB40 = R9C20_GBO1;
assign R2C23_GB40 = R2C24_GBO1;
assign R2C24_GB40 = R2C24_GBO1;
assign R2C25_GB40 = R2C24_GBO1;
assign R2C26_GB40 = R2C24_GBO1;
assign R2C27_GB40 = R2C24_GBO1;
assign R2C28_GB40 = R2C24_GBO1;
assign R3C23_GB40 = R3C24_GBO1;
assign R3C24_GB40 = R3C24_GBO1;
assign R3C25_GB40 = R3C24_GBO1;
assign R3C26_GB40 = R3C24_GBO1;
assign R3C27_GB40 = R3C24_GBO1;
assign R3C28_GB40 = R3C24_GBO1;
assign R4C23_GB40 = R4C24_GBO1;
assign R4C24_GB40 = R4C24_GBO1;
assign R4C25_GB40 = R4C24_GBO1;
assign R4C26_GB40 = R4C24_GBO1;
assign R4C27_GB40 = R4C24_GBO1;
assign R4C28_GB40 = R4C24_GBO1;
assign R5C23_GB40 = R5C24_GBO1;
assign R5C24_GB40 = R5C24_GBO1;
assign R5C25_GB40 = R5C24_GBO1;
assign R5C26_GB40 = R5C24_GBO1;
assign R5C27_GB40 = R5C24_GBO1;
assign R5C28_GB40 = R5C24_GBO1;
assign R6C23_GB40 = R6C24_GBO1;
assign R6C24_GB40 = R6C24_GBO1;
assign R6C25_GB40 = R6C24_GBO1;
assign R6C26_GB40 = R6C24_GBO1;
assign R6C27_GB40 = R6C24_GBO1;
assign R6C28_GB40 = R6C24_GBO1;
assign R7C23_GB40 = R7C24_GBO1;
assign R7C24_GB40 = R7C24_GBO1;
assign R7C25_GB40 = R7C24_GBO1;
assign R7C26_GB40 = R7C24_GBO1;
assign R7C27_GB40 = R7C24_GBO1;
assign R7C28_GB40 = R7C24_GBO1;
assign R8C23_GB40 = R8C24_GBO1;
assign R8C24_GB40 = R8C24_GBO1;
assign R8C25_GB40 = R8C24_GBO1;
assign R8C26_GB40 = R8C24_GBO1;
assign R8C27_GB40 = R8C24_GBO1;
assign R8C28_GB40 = R8C24_GBO1;
assign R9C23_GB40 = R9C24_GBO1;
assign R9C24_GB40 = R9C24_GBO1;
assign R9C25_GB40 = R9C24_GBO1;
assign R9C26_GB40 = R9C24_GBO1;
assign R9C27_GB40 = R9C24_GBO1;
assign R9C28_GB40 = R9C24_GBO1;
assign R2C2_GB50 = R2C3_GBO1;
assign R2C3_GB50 = R2C3_GBO1;
assign R2C4_GB50 = R2C3_GBO1;
assign R2C5_GB50 = R2C3_GBO1;
assign R3C2_GB50 = R3C3_GBO1;
assign R3C3_GB50 = R3C3_GBO1;
assign R3C4_GB50 = R3C3_GBO1;
assign R3C5_GB50 = R3C3_GBO1;
assign R4C2_GB50 = R4C3_GBO1;
assign R4C3_GB50 = R4C3_GBO1;
assign R4C4_GB50 = R4C3_GBO1;
assign R4C5_GB50 = R4C3_GBO1;
assign R5C2_GB50 = R5C3_GBO1;
assign R5C3_GB50 = R5C3_GBO1;
assign R5C4_GB50 = R5C3_GBO1;
assign R5C5_GB50 = R5C3_GBO1;
assign R6C2_GB50 = R6C3_GBO1;
assign R6C3_GB50 = R6C3_GBO1;
assign R6C4_GB50 = R6C3_GBO1;
assign R6C5_GB50 = R6C3_GBO1;
assign R7C2_GB50 = R7C3_GBO1;
assign R7C3_GB50 = R7C3_GBO1;
assign R7C4_GB50 = R7C3_GBO1;
assign R7C5_GB50 = R7C3_GBO1;
assign R8C2_GB50 = R8C3_GBO1;
assign R8C3_GB50 = R8C3_GBO1;
assign R8C4_GB50 = R8C3_GBO1;
assign R8C5_GB50 = R8C3_GBO1;
assign R9C2_GB50 = R9C3_GBO1;
assign R9C3_GB50 = R9C3_GBO1;
assign R9C4_GB50 = R9C3_GBO1;
assign R9C5_GB50 = R9C3_GBO1;
assign R2C9_GB50 = R2C7_GBO1;
assign R2C6_GB50 = R2C7_GBO1;
assign R2C7_GB50 = R2C7_GBO1;
assign R2C8_GB50 = R2C7_GBO1;
assign R3C9_GB50 = R3C7_GBO1;
assign R3C6_GB50 = R3C7_GBO1;
assign R3C7_GB50 = R3C7_GBO1;
assign R3C8_GB50 = R3C7_GBO1;
assign R4C9_GB50 = R4C7_GBO1;
assign R4C6_GB50 = R4C7_GBO1;
assign R4C7_GB50 = R4C7_GBO1;
assign R4C8_GB50 = R4C7_GBO1;
assign R5C9_GB50 = R5C7_GBO1;
assign R5C6_GB50 = R5C7_GBO1;
assign R5C7_GB50 = R5C7_GBO1;
assign R5C8_GB50 = R5C7_GBO1;
assign R6C9_GB50 = R6C7_GBO1;
assign R6C6_GB50 = R6C7_GBO1;
assign R6C7_GB50 = R6C7_GBO1;
assign R6C8_GB50 = R6C7_GBO1;
assign R7C9_GB50 = R7C7_GBO1;
assign R7C6_GB50 = R7C7_GBO1;
assign R7C7_GB50 = R7C7_GBO1;
assign R7C8_GB50 = R7C7_GBO1;
assign R8C9_GB50 = R8C7_GBO1;
assign R8C6_GB50 = R8C7_GBO1;
assign R8C7_GB50 = R8C7_GBO1;
assign R8C8_GB50 = R8C7_GBO1;
assign R9C9_GB50 = R9C7_GBO1;
assign R9C6_GB50 = R9C7_GBO1;
assign R9C7_GB50 = R9C7_GBO1;
assign R9C8_GB50 = R9C7_GBO1;
assign R2C10_GB50 = R2C11_GBO1;
assign R2C11_GB50 = R2C11_GBO1;
assign R2C12_GB50 = R2C11_GBO1;
assign R2C13_GB50 = R2C11_GBO1;
assign R3C10_GB50 = R3C11_GBO1;
assign R3C11_GB50 = R3C11_GBO1;
assign R3C12_GB50 = R3C11_GBO1;
assign R3C13_GB50 = R3C11_GBO1;
assign R4C10_GB50 = R4C11_GBO1;
assign R4C11_GB50 = R4C11_GBO1;
assign R4C12_GB50 = R4C11_GBO1;
assign R4C13_GB50 = R4C11_GBO1;
assign R5C10_GB50 = R5C11_GBO1;
assign R5C11_GB50 = R5C11_GBO1;
assign R5C12_GB50 = R5C11_GBO1;
assign R5C13_GB50 = R5C11_GBO1;
assign R6C10_GB50 = R6C11_GBO1;
assign R6C11_GB50 = R6C11_GBO1;
assign R6C12_GB50 = R6C11_GBO1;
assign R6C13_GB50 = R6C11_GBO1;
assign R7C10_GB50 = R7C11_GBO1;
assign R7C11_GB50 = R7C11_GBO1;
assign R7C12_GB50 = R7C11_GBO1;
assign R7C13_GB50 = R7C11_GBO1;
assign R8C10_GB50 = R8C11_GBO1;
assign R8C11_GB50 = R8C11_GBO1;
assign R8C12_GB50 = R8C11_GBO1;
assign R8C13_GB50 = R8C11_GBO1;
assign R9C10_GB50 = R9C11_GBO1;
assign R9C11_GB50 = R9C11_GBO1;
assign R9C12_GB50 = R9C11_GBO1;
assign R9C13_GB50 = R9C11_GBO1;
assign R2C17_GB50 = R2C15_GBO1;
assign R2C14_GB50 = R2C15_GBO1;
assign R2C15_GB50 = R2C15_GBO1;
assign R2C16_GB50 = R2C15_GBO1;
assign R3C17_GB50 = R3C15_GBO1;
assign R3C14_GB50 = R3C15_GBO1;
assign R3C15_GB50 = R3C15_GBO1;
assign R3C16_GB50 = R3C15_GBO1;
assign R4C17_GB50 = R4C15_GBO1;
assign R4C14_GB50 = R4C15_GBO1;
assign R4C15_GB50 = R4C15_GBO1;
assign R4C16_GB50 = R4C15_GBO1;
assign R5C17_GB50 = R5C15_GBO1;
assign R5C14_GB50 = R5C15_GBO1;
assign R5C15_GB50 = R5C15_GBO1;
assign R5C16_GB50 = R5C15_GBO1;
assign R6C17_GB50 = R6C15_GBO1;
assign R6C14_GB50 = R6C15_GBO1;
assign R6C15_GB50 = R6C15_GBO1;
assign R6C16_GB50 = R6C15_GBO1;
assign R7C17_GB50 = R7C15_GBO1;
assign R7C14_GB50 = R7C15_GBO1;
assign R7C15_GB50 = R7C15_GBO1;
assign R7C16_GB50 = R7C15_GBO1;
assign R8C17_GB50 = R8C15_GBO1;
assign R8C14_GB50 = R8C15_GBO1;
assign R8C15_GB50 = R8C15_GBO1;
assign R8C16_GB50 = R8C15_GBO1;
assign R9C17_GB50 = R9C15_GBO1;
assign R9C14_GB50 = R9C15_GBO1;
assign R9C15_GB50 = R9C15_GBO1;
assign R9C16_GB50 = R9C15_GBO1;
assign R2C18_GB50 = R2C19_GBO1;
assign R2C19_GB50 = R2C19_GBO1;
assign R2C20_GB50 = R2C19_GBO1;
assign R2C21_GB50 = R2C19_GBO1;
assign R3C18_GB50 = R3C19_GBO1;
assign R3C19_GB50 = R3C19_GBO1;
assign R3C20_GB50 = R3C19_GBO1;
assign R3C21_GB50 = R3C19_GBO1;
assign R4C18_GB50 = R4C19_GBO1;
assign R4C19_GB50 = R4C19_GBO1;
assign R4C20_GB50 = R4C19_GBO1;
assign R4C21_GB50 = R4C19_GBO1;
assign R5C18_GB50 = R5C19_GBO1;
assign R5C19_GB50 = R5C19_GBO1;
assign R5C20_GB50 = R5C19_GBO1;
assign R5C21_GB50 = R5C19_GBO1;
assign R6C18_GB50 = R6C19_GBO1;
assign R6C19_GB50 = R6C19_GBO1;
assign R6C20_GB50 = R6C19_GBO1;
assign R6C21_GB50 = R6C19_GBO1;
assign R7C18_GB50 = R7C19_GBO1;
assign R7C19_GB50 = R7C19_GBO1;
assign R7C20_GB50 = R7C19_GBO1;
assign R7C21_GB50 = R7C19_GBO1;
assign R8C18_GB50 = R8C19_GBO1;
assign R8C19_GB50 = R8C19_GBO1;
assign R8C20_GB50 = R8C19_GBO1;
assign R8C21_GB50 = R8C19_GBO1;
assign R9C18_GB50 = R9C19_GBO1;
assign R9C19_GB50 = R9C19_GBO1;
assign R9C20_GB50 = R9C19_GBO1;
assign R9C21_GB50 = R9C19_GBO1;
assign R2C25_GB50 = R2C23_GBO1;
assign R2C22_GB50 = R2C23_GBO1;
assign R2C23_GB50 = R2C23_GBO1;
assign R2C24_GB50 = R2C23_GBO1;
assign R3C25_GB50 = R3C23_GBO1;
assign R3C22_GB50 = R3C23_GBO1;
assign R3C23_GB50 = R3C23_GBO1;
assign R3C24_GB50 = R3C23_GBO1;
assign R4C25_GB50 = R4C23_GBO1;
assign R4C22_GB50 = R4C23_GBO1;
assign R4C23_GB50 = R4C23_GBO1;
assign R4C24_GB50 = R4C23_GBO1;
assign R5C25_GB50 = R5C23_GBO1;
assign R5C22_GB50 = R5C23_GBO1;
assign R5C23_GB50 = R5C23_GBO1;
assign R5C24_GB50 = R5C23_GBO1;
assign R6C25_GB50 = R6C23_GBO1;
assign R6C22_GB50 = R6C23_GBO1;
assign R6C23_GB50 = R6C23_GBO1;
assign R6C24_GB50 = R6C23_GBO1;
assign R7C25_GB50 = R7C23_GBO1;
assign R7C22_GB50 = R7C23_GBO1;
assign R7C23_GB50 = R7C23_GBO1;
assign R7C24_GB50 = R7C23_GBO1;
assign R8C25_GB50 = R8C23_GBO1;
assign R8C22_GB50 = R8C23_GBO1;
assign R8C23_GB50 = R8C23_GBO1;
assign R8C24_GB50 = R8C23_GBO1;
assign R9C25_GB50 = R9C23_GBO1;
assign R9C22_GB50 = R9C23_GBO1;
assign R9C23_GB50 = R9C23_GBO1;
assign R9C24_GB50 = R9C23_GBO1;
assign R2C26_GB50 = R2C27_GBO1;
assign R2C27_GB50 = R2C27_GBO1;
assign R2C28_GB50 = R2C27_GBO1;
assign R3C26_GB50 = R3C27_GBO1;
assign R3C27_GB50 = R3C27_GBO1;
assign R3C28_GB50 = R3C27_GBO1;
assign R4C26_GB50 = R4C27_GBO1;
assign R4C27_GB50 = R4C27_GBO1;
assign R4C28_GB50 = R4C27_GBO1;
assign R5C26_GB50 = R5C27_GBO1;
assign R5C27_GB50 = R5C27_GBO1;
assign R5C28_GB50 = R5C27_GBO1;
assign R6C26_GB50 = R6C27_GBO1;
assign R6C27_GB50 = R6C27_GBO1;
assign R6C28_GB50 = R6C27_GBO1;
assign R7C26_GB50 = R7C27_GBO1;
assign R7C27_GB50 = R7C27_GBO1;
assign R7C28_GB50 = R7C27_GBO1;
assign R8C26_GB50 = R8C27_GBO1;
assign R8C27_GB50 = R8C27_GBO1;
assign R8C28_GB50 = R8C27_GBO1;
assign R9C26_GB50 = R9C27_GBO1;
assign R9C27_GB50 = R9C27_GBO1;
assign R9C28_GB50 = R9C27_GBO1;
assign R2C2_GB60 = R2C2_GBO1;
assign R2C3_GB60 = R2C2_GBO1;
assign R2C4_GB60 = R2C2_GBO1;
assign R3C2_GB60 = R3C2_GBO1;
assign R3C3_GB60 = R3C2_GBO1;
assign R3C4_GB60 = R3C2_GBO1;
assign R4C2_GB60 = R4C2_GBO1;
assign R4C3_GB60 = R4C2_GBO1;
assign R4C4_GB60 = R4C2_GBO1;
assign R5C2_GB60 = R5C2_GBO1;
assign R5C3_GB60 = R5C2_GBO1;
assign R5C4_GB60 = R5C2_GBO1;
assign R6C2_GB60 = R6C2_GBO1;
assign R6C3_GB60 = R6C2_GBO1;
assign R6C4_GB60 = R6C2_GBO1;
assign R7C2_GB60 = R7C2_GBO1;
assign R7C3_GB60 = R7C2_GBO1;
assign R7C4_GB60 = R7C2_GBO1;
assign R8C2_GB60 = R8C2_GBO1;
assign R8C3_GB60 = R8C2_GBO1;
assign R8C4_GB60 = R8C2_GBO1;
assign R9C2_GB60 = R9C2_GBO1;
assign R9C3_GB60 = R9C2_GBO1;
assign R9C4_GB60 = R9C2_GBO1;
assign R2C5_GB60 = R2C6_GBO1;
assign R2C6_GB60 = R2C6_GBO1;
assign R2C7_GB60 = R2C6_GBO1;
assign R2C8_GB60 = R2C6_GBO1;
assign R3C5_GB60 = R3C6_GBO1;
assign R3C6_GB60 = R3C6_GBO1;
assign R3C7_GB60 = R3C6_GBO1;
assign R3C8_GB60 = R3C6_GBO1;
assign R4C5_GB60 = R4C6_GBO1;
assign R4C6_GB60 = R4C6_GBO1;
assign R4C7_GB60 = R4C6_GBO1;
assign R4C8_GB60 = R4C6_GBO1;
assign R5C5_GB60 = R5C6_GBO1;
assign R5C6_GB60 = R5C6_GBO1;
assign R5C7_GB60 = R5C6_GBO1;
assign R5C8_GB60 = R5C6_GBO1;
assign R6C5_GB60 = R6C6_GBO1;
assign R6C6_GB60 = R6C6_GBO1;
assign R6C7_GB60 = R6C6_GBO1;
assign R6C8_GB60 = R6C6_GBO1;
assign R7C5_GB60 = R7C6_GBO1;
assign R7C6_GB60 = R7C6_GBO1;
assign R7C7_GB60 = R7C6_GBO1;
assign R7C8_GB60 = R7C6_GBO1;
assign R8C5_GB60 = R8C6_GBO1;
assign R8C6_GB60 = R8C6_GBO1;
assign R8C7_GB60 = R8C6_GBO1;
assign R8C8_GB60 = R8C6_GBO1;
assign R9C5_GB60 = R9C6_GBO1;
assign R9C6_GB60 = R9C6_GBO1;
assign R9C7_GB60 = R9C6_GBO1;
assign R9C8_GB60 = R9C6_GBO1;
assign R2C9_GB60 = R2C10_GBO1;
assign R2C10_GB60 = R2C10_GBO1;
assign R2C11_GB60 = R2C10_GBO1;
assign R2C12_GB60 = R2C10_GBO1;
assign R3C9_GB60 = R3C10_GBO1;
assign R3C10_GB60 = R3C10_GBO1;
assign R3C11_GB60 = R3C10_GBO1;
assign R3C12_GB60 = R3C10_GBO1;
assign R4C9_GB60 = R4C10_GBO1;
assign R4C10_GB60 = R4C10_GBO1;
assign R4C11_GB60 = R4C10_GBO1;
assign R4C12_GB60 = R4C10_GBO1;
assign R5C9_GB60 = R5C10_GBO1;
assign R5C10_GB60 = R5C10_GBO1;
assign R5C11_GB60 = R5C10_GBO1;
assign R5C12_GB60 = R5C10_GBO1;
assign R6C9_GB60 = R6C10_GBO1;
assign R6C10_GB60 = R6C10_GBO1;
assign R6C11_GB60 = R6C10_GBO1;
assign R6C12_GB60 = R6C10_GBO1;
assign R7C9_GB60 = R7C10_GBO1;
assign R7C10_GB60 = R7C10_GBO1;
assign R7C11_GB60 = R7C10_GBO1;
assign R7C12_GB60 = R7C10_GBO1;
assign R8C9_GB60 = R8C10_GBO1;
assign R8C10_GB60 = R8C10_GBO1;
assign R8C11_GB60 = R8C10_GBO1;
assign R8C12_GB60 = R8C10_GBO1;
assign R9C9_GB60 = R9C10_GBO1;
assign R9C10_GB60 = R9C10_GBO1;
assign R9C11_GB60 = R9C10_GBO1;
assign R9C12_GB60 = R9C10_GBO1;
assign R2C13_GB60 = R2C14_GBO1;
assign R2C14_GB60 = R2C14_GBO1;
assign R2C15_GB60 = R2C14_GBO1;
assign R2C16_GB60 = R2C14_GBO1;
assign R3C13_GB60 = R3C14_GBO1;
assign R3C14_GB60 = R3C14_GBO1;
assign R3C15_GB60 = R3C14_GBO1;
assign R3C16_GB60 = R3C14_GBO1;
assign R4C13_GB60 = R4C14_GBO1;
assign R4C14_GB60 = R4C14_GBO1;
assign R4C15_GB60 = R4C14_GBO1;
assign R4C16_GB60 = R4C14_GBO1;
assign R5C13_GB60 = R5C14_GBO1;
assign R5C14_GB60 = R5C14_GBO1;
assign R5C15_GB60 = R5C14_GBO1;
assign R5C16_GB60 = R5C14_GBO1;
assign R6C13_GB60 = R6C14_GBO1;
assign R6C14_GB60 = R6C14_GBO1;
assign R6C15_GB60 = R6C14_GBO1;
assign R6C16_GB60 = R6C14_GBO1;
assign R7C13_GB60 = R7C14_GBO1;
assign R7C14_GB60 = R7C14_GBO1;
assign R7C15_GB60 = R7C14_GBO1;
assign R7C16_GB60 = R7C14_GBO1;
assign R8C13_GB60 = R8C14_GBO1;
assign R8C14_GB60 = R8C14_GBO1;
assign R8C15_GB60 = R8C14_GBO1;
assign R8C16_GB60 = R8C14_GBO1;
assign R9C13_GB60 = R9C14_GBO1;
assign R9C14_GB60 = R9C14_GBO1;
assign R9C15_GB60 = R9C14_GBO1;
assign R9C16_GB60 = R9C14_GBO1;
assign R2C17_GB60 = R2C18_GBO1;
assign R2C18_GB60 = R2C18_GBO1;
assign R2C19_GB60 = R2C18_GBO1;
assign R2C20_GB60 = R2C18_GBO1;
assign R3C17_GB60 = R3C18_GBO1;
assign R3C18_GB60 = R3C18_GBO1;
assign R3C19_GB60 = R3C18_GBO1;
assign R3C20_GB60 = R3C18_GBO1;
assign R4C17_GB60 = R4C18_GBO1;
assign R4C18_GB60 = R4C18_GBO1;
assign R4C19_GB60 = R4C18_GBO1;
assign R4C20_GB60 = R4C18_GBO1;
assign R5C17_GB60 = R5C18_GBO1;
assign R5C18_GB60 = R5C18_GBO1;
assign R5C19_GB60 = R5C18_GBO1;
assign R5C20_GB60 = R5C18_GBO1;
assign R6C17_GB60 = R6C18_GBO1;
assign R6C18_GB60 = R6C18_GBO1;
assign R6C19_GB60 = R6C18_GBO1;
assign R6C20_GB60 = R6C18_GBO1;
assign R7C17_GB60 = R7C18_GBO1;
assign R7C18_GB60 = R7C18_GBO1;
assign R7C19_GB60 = R7C18_GBO1;
assign R7C20_GB60 = R7C18_GBO1;
assign R8C17_GB60 = R8C18_GBO1;
assign R8C18_GB60 = R8C18_GBO1;
assign R8C19_GB60 = R8C18_GBO1;
assign R8C20_GB60 = R8C18_GBO1;
assign R9C17_GB60 = R9C18_GBO1;
assign R9C18_GB60 = R9C18_GBO1;
assign R9C19_GB60 = R9C18_GBO1;
assign R9C20_GB60 = R9C18_GBO1;
assign R2C21_GB60 = R2C22_GBO1;
assign R2C22_GB60 = R2C22_GBO1;
assign R2C23_GB60 = R2C22_GBO1;
assign R2C24_GB60 = R2C22_GBO1;
assign R3C21_GB60 = R3C22_GBO1;
assign R3C22_GB60 = R3C22_GBO1;
assign R3C23_GB60 = R3C22_GBO1;
assign R3C24_GB60 = R3C22_GBO1;
assign R4C21_GB60 = R4C22_GBO1;
assign R4C22_GB60 = R4C22_GBO1;
assign R4C23_GB60 = R4C22_GBO1;
assign R4C24_GB60 = R4C22_GBO1;
assign R5C21_GB60 = R5C22_GBO1;
assign R5C22_GB60 = R5C22_GBO1;
assign R5C23_GB60 = R5C22_GBO1;
assign R5C24_GB60 = R5C22_GBO1;
assign R6C21_GB60 = R6C22_GBO1;
assign R6C22_GB60 = R6C22_GBO1;
assign R6C23_GB60 = R6C22_GBO1;
assign R6C24_GB60 = R6C22_GBO1;
assign R7C21_GB60 = R7C22_GBO1;
assign R7C22_GB60 = R7C22_GBO1;
assign R7C23_GB60 = R7C22_GBO1;
assign R7C24_GB60 = R7C22_GBO1;
assign R8C21_GB60 = R8C22_GBO1;
assign R8C22_GB60 = R8C22_GBO1;
assign R8C23_GB60 = R8C22_GBO1;
assign R8C24_GB60 = R8C22_GBO1;
assign R9C21_GB60 = R9C22_GBO1;
assign R9C22_GB60 = R9C22_GBO1;
assign R9C23_GB60 = R9C22_GBO1;
assign R9C24_GB60 = R9C22_GBO1;
assign R2C25_GB60 = R2C26_GBO1;
assign R2C26_GB60 = R2C26_GBO1;
assign R2C27_GB60 = R2C26_GBO1;
assign R2C28_GB60 = R2C26_GBO1;
assign R3C25_GB60 = R3C26_GBO1;
assign R3C26_GB60 = R3C26_GBO1;
assign R3C27_GB60 = R3C26_GBO1;
assign R3C28_GB60 = R3C26_GBO1;
assign R4C25_GB60 = R4C26_GBO1;
assign R4C26_GB60 = R4C26_GBO1;
assign R4C27_GB60 = R4C26_GBO1;
assign R4C28_GB60 = R4C26_GBO1;
assign R5C25_GB60 = R5C26_GBO1;
assign R5C26_GB60 = R5C26_GBO1;
assign R5C27_GB60 = R5C26_GBO1;
assign R5C28_GB60 = R5C26_GBO1;
assign R6C25_GB60 = R6C26_GBO1;
assign R6C26_GB60 = R6C26_GBO1;
assign R6C27_GB60 = R6C26_GBO1;
assign R6C28_GB60 = R6C26_GBO1;
assign R7C25_GB60 = R7C26_GBO1;
assign R7C26_GB60 = R7C26_GBO1;
assign R7C27_GB60 = R7C26_GBO1;
assign R7C28_GB60 = R7C26_GBO1;
assign R8C25_GB60 = R8C26_GBO1;
assign R8C26_GB60 = R8C26_GBO1;
assign R8C27_GB60 = R8C26_GBO1;
assign R8C28_GB60 = R8C26_GBO1;
assign R9C25_GB60 = R9C26_GBO1;
assign R9C26_GB60 = R9C26_GBO1;
assign R9C27_GB60 = R9C26_GBO1;
assign R9C28_GB60 = R9C26_GBO1;
assign R2C2_GB70 = R2C1_GBO1;
assign R2C3_GB70 = R2C1_GBO1;
assign R3C2_GB70 = R3C1_GBO1;
assign R3C3_GB70 = R3C1_GBO1;
assign R4C2_GB70 = R4C1_GBO1;
assign R4C3_GB70 = R4C1_GBO1;
assign R5C2_GB70 = R5C1_GBO1;
assign R5C3_GB70 = R5C1_GBO1;
assign R6C2_GB70 = R6C1_GBO1;
assign R6C3_GB70 = R6C1_GBO1;
assign R7C2_GB70 = R7C1_GBO1;
assign R7C3_GB70 = R7C1_GBO1;
assign R8C2_GB70 = R8C1_GBO1;
assign R8C3_GB70 = R8C1_GBO1;
assign R9C2_GB70 = R9C1_GBO1;
assign R9C3_GB70 = R9C1_GBO1;
assign R2C4_GB70 = R2C5_GBO1;
assign R2C5_GB70 = R2C5_GBO1;
assign R2C6_GB70 = R2C5_GBO1;
assign R2C7_GB70 = R2C5_GBO1;
assign R3C4_GB70 = R3C5_GBO1;
assign R3C5_GB70 = R3C5_GBO1;
assign R3C6_GB70 = R3C5_GBO1;
assign R3C7_GB70 = R3C5_GBO1;
assign R4C4_GB70 = R4C5_GBO1;
assign R4C5_GB70 = R4C5_GBO1;
assign R4C6_GB70 = R4C5_GBO1;
assign R4C7_GB70 = R4C5_GBO1;
assign R5C4_GB70 = R5C5_GBO1;
assign R5C5_GB70 = R5C5_GBO1;
assign R5C6_GB70 = R5C5_GBO1;
assign R5C7_GB70 = R5C5_GBO1;
assign R6C4_GB70 = R6C5_GBO1;
assign R6C5_GB70 = R6C5_GBO1;
assign R6C6_GB70 = R6C5_GBO1;
assign R6C7_GB70 = R6C5_GBO1;
assign R7C4_GB70 = R7C5_GBO1;
assign R7C5_GB70 = R7C5_GBO1;
assign R7C6_GB70 = R7C5_GBO1;
assign R7C7_GB70 = R7C5_GBO1;
assign R8C4_GB70 = R8C5_GBO1;
assign R8C5_GB70 = R8C5_GBO1;
assign R8C6_GB70 = R8C5_GBO1;
assign R8C7_GB70 = R8C5_GBO1;
assign R9C4_GB70 = R9C5_GBO1;
assign R9C5_GB70 = R9C5_GBO1;
assign R9C6_GB70 = R9C5_GBO1;
assign R9C7_GB70 = R9C5_GBO1;
assign R2C9_GB70 = R2C9_GBO1;
assign R2C10_GB70 = R2C9_GBO1;
assign R2C11_GB70 = R2C9_GBO1;
assign R2C8_GB70 = R2C9_GBO1;
assign R3C9_GB70 = R3C9_GBO1;
assign R3C10_GB70 = R3C9_GBO1;
assign R3C11_GB70 = R3C9_GBO1;
assign R3C8_GB70 = R3C9_GBO1;
assign R4C9_GB70 = R4C9_GBO1;
assign R4C10_GB70 = R4C9_GBO1;
assign R4C11_GB70 = R4C9_GBO1;
assign R4C8_GB70 = R4C9_GBO1;
assign R5C9_GB70 = R5C9_GBO1;
assign R5C10_GB70 = R5C9_GBO1;
assign R5C11_GB70 = R5C9_GBO1;
assign R5C8_GB70 = R5C9_GBO1;
assign R6C9_GB70 = R6C9_GBO1;
assign R6C10_GB70 = R6C9_GBO1;
assign R6C11_GB70 = R6C9_GBO1;
assign R6C8_GB70 = R6C9_GBO1;
assign R7C9_GB70 = R7C9_GBO1;
assign R7C10_GB70 = R7C9_GBO1;
assign R7C11_GB70 = R7C9_GBO1;
assign R7C8_GB70 = R7C9_GBO1;
assign R8C9_GB70 = R8C9_GBO1;
assign R8C10_GB70 = R8C9_GBO1;
assign R8C11_GB70 = R8C9_GBO1;
assign R8C8_GB70 = R8C9_GBO1;
assign R9C9_GB70 = R9C9_GBO1;
assign R9C10_GB70 = R9C9_GBO1;
assign R9C11_GB70 = R9C9_GBO1;
assign R9C8_GB70 = R9C9_GBO1;
assign R2C12_GB70 = R2C13_GBO1;
assign R2C13_GB70 = R2C13_GBO1;
assign R2C14_GB70 = R2C13_GBO1;
assign R2C15_GB70 = R2C13_GBO1;
assign R3C12_GB70 = R3C13_GBO1;
assign R3C13_GB70 = R3C13_GBO1;
assign R3C14_GB70 = R3C13_GBO1;
assign R3C15_GB70 = R3C13_GBO1;
assign R4C12_GB70 = R4C13_GBO1;
assign R4C13_GB70 = R4C13_GBO1;
assign R4C14_GB70 = R4C13_GBO1;
assign R4C15_GB70 = R4C13_GBO1;
assign R5C12_GB70 = R5C13_GBO1;
assign R5C13_GB70 = R5C13_GBO1;
assign R5C14_GB70 = R5C13_GBO1;
assign R5C15_GB70 = R5C13_GBO1;
assign R6C12_GB70 = R6C13_GBO1;
assign R6C13_GB70 = R6C13_GBO1;
assign R6C14_GB70 = R6C13_GBO1;
assign R6C15_GB70 = R6C13_GBO1;
assign R7C12_GB70 = R7C13_GBO1;
assign R7C13_GB70 = R7C13_GBO1;
assign R7C14_GB70 = R7C13_GBO1;
assign R7C15_GB70 = R7C13_GBO1;
assign R8C12_GB70 = R8C13_GBO1;
assign R8C13_GB70 = R8C13_GBO1;
assign R8C14_GB70 = R8C13_GBO1;
assign R8C15_GB70 = R8C13_GBO1;
assign R9C12_GB70 = R9C13_GBO1;
assign R9C13_GB70 = R9C13_GBO1;
assign R9C14_GB70 = R9C13_GBO1;
assign R9C15_GB70 = R9C13_GBO1;
assign R2C17_GB70 = R2C17_GBO1;
assign R2C18_GB70 = R2C17_GBO1;
assign R2C19_GB70 = R2C17_GBO1;
assign R2C16_GB70 = R2C17_GBO1;
assign R3C17_GB70 = R3C17_GBO1;
assign R3C18_GB70 = R3C17_GBO1;
assign R3C19_GB70 = R3C17_GBO1;
assign R3C16_GB70 = R3C17_GBO1;
assign R4C17_GB70 = R4C17_GBO1;
assign R4C18_GB70 = R4C17_GBO1;
assign R4C19_GB70 = R4C17_GBO1;
assign R4C16_GB70 = R4C17_GBO1;
assign R5C17_GB70 = R5C17_GBO1;
assign R5C18_GB70 = R5C17_GBO1;
assign R5C19_GB70 = R5C17_GBO1;
assign R5C16_GB70 = R5C17_GBO1;
assign R6C17_GB70 = R6C17_GBO1;
assign R6C18_GB70 = R6C17_GBO1;
assign R6C19_GB70 = R6C17_GBO1;
assign R6C16_GB70 = R6C17_GBO1;
assign R7C17_GB70 = R7C17_GBO1;
assign R7C18_GB70 = R7C17_GBO1;
assign R7C19_GB70 = R7C17_GBO1;
assign R7C16_GB70 = R7C17_GBO1;
assign R8C17_GB70 = R8C17_GBO1;
assign R8C18_GB70 = R8C17_GBO1;
assign R8C19_GB70 = R8C17_GBO1;
assign R8C16_GB70 = R8C17_GBO1;
assign R9C17_GB70 = R9C17_GBO1;
assign R9C18_GB70 = R9C17_GBO1;
assign R9C19_GB70 = R9C17_GBO1;
assign R9C16_GB70 = R9C17_GBO1;
assign R2C20_GB70 = R2C21_GBO1;
assign R2C21_GB70 = R2C21_GBO1;
assign R2C22_GB70 = R2C21_GBO1;
assign R2C23_GB70 = R2C21_GBO1;
assign R3C20_GB70 = R3C21_GBO1;
assign R3C21_GB70 = R3C21_GBO1;
assign R3C22_GB70 = R3C21_GBO1;
assign R3C23_GB70 = R3C21_GBO1;
assign R4C20_GB70 = R4C21_GBO1;
assign R4C21_GB70 = R4C21_GBO1;
assign R4C22_GB70 = R4C21_GBO1;
assign R4C23_GB70 = R4C21_GBO1;
assign R5C20_GB70 = R5C21_GBO1;
assign R5C21_GB70 = R5C21_GBO1;
assign R5C22_GB70 = R5C21_GBO1;
assign R5C23_GB70 = R5C21_GBO1;
assign R6C20_GB70 = R6C21_GBO1;
assign R6C21_GB70 = R6C21_GBO1;
assign R6C22_GB70 = R6C21_GBO1;
assign R6C23_GB70 = R6C21_GBO1;
assign R7C20_GB70 = R7C21_GBO1;
assign R7C21_GB70 = R7C21_GBO1;
assign R7C22_GB70 = R7C21_GBO1;
assign R7C23_GB70 = R7C21_GBO1;
assign R8C20_GB70 = R8C21_GBO1;
assign R8C21_GB70 = R8C21_GBO1;
assign R8C22_GB70 = R8C21_GBO1;
assign R8C23_GB70 = R8C21_GBO1;
assign R9C20_GB70 = R9C21_GBO1;
assign R9C21_GB70 = R9C21_GBO1;
assign R9C22_GB70 = R9C21_GBO1;
assign R9C23_GB70 = R9C21_GBO1;
assign R2C24_GB70 = R2C25_GBO1;
assign R2C25_GB70 = R2C25_GBO1;
assign R2C26_GB70 = R2C25_GBO1;
assign R2C27_GB70 = R2C25_GBO1;
assign R2C28_GB70 = R2C25_GBO1;
assign R3C24_GB70 = R3C25_GBO1;
assign R3C25_GB70 = R3C25_GBO1;
assign R3C26_GB70 = R3C25_GBO1;
assign R3C27_GB70 = R3C25_GBO1;
assign R3C28_GB70 = R3C25_GBO1;
assign R4C24_GB70 = R4C25_GBO1;
assign R4C25_GB70 = R4C25_GBO1;
assign R4C26_GB70 = R4C25_GBO1;
assign R4C27_GB70 = R4C25_GBO1;
assign R4C28_GB70 = R4C25_GBO1;
assign R5C24_GB70 = R5C25_GBO1;
assign R5C25_GB70 = R5C25_GBO1;
assign R5C26_GB70 = R5C25_GBO1;
assign R5C27_GB70 = R5C25_GBO1;
assign R5C28_GB70 = R5C25_GBO1;
assign R6C24_GB70 = R6C25_GBO1;
assign R6C25_GB70 = R6C25_GBO1;
assign R6C26_GB70 = R6C25_GBO1;
assign R6C27_GB70 = R6C25_GBO1;
assign R6C28_GB70 = R6C25_GBO1;
assign R7C24_GB70 = R7C25_GBO1;
assign R7C25_GB70 = R7C25_GBO1;
assign R7C26_GB70 = R7C25_GBO1;
assign R7C27_GB70 = R7C25_GBO1;
assign R7C28_GB70 = R7C25_GBO1;
assign R8C24_GB70 = R8C25_GBO1;
assign R8C25_GB70 = R8C25_GBO1;
assign R8C26_GB70 = R8C25_GBO1;
assign R8C27_GB70 = R8C25_GBO1;
assign R8C28_GB70 = R8C25_GBO1;
assign R9C24_GB70 = R9C25_GBO1;
assign R9C25_GB70 = R9C25_GBO1;
assign R9C26_GB70 = R9C25_GBO1;
assign R9C27_GB70 = R9C25_GBO1;
assign R9C28_GB70 = R9C25_GBO1;
assign R11C2_GB00 = R11C4_GBO0;
assign R11C3_GB00 = R11C4_GBO0;
assign R11C4_GB00 = R11C4_GBO0;
assign R11C5_GB00 = R11C4_GBO0;
assign R11C6_GB00 = R11C4_GBO0;
assign R12C2_GB00 = R12C4_GBO0;
assign R12C3_GB00 = R12C4_GBO0;
assign R12C4_GB00 = R12C4_GBO0;
assign R12C5_GB00 = R12C4_GBO0;
assign R12C6_GB00 = R12C4_GBO0;
assign R13C2_GB00 = R13C4_GBO0;
assign R13C3_GB00 = R13C4_GBO0;
assign R13C4_GB00 = R13C4_GBO0;
assign R13C5_GB00 = R13C4_GBO0;
assign R13C6_GB00 = R13C4_GBO0;
assign R14C2_GB00 = R14C4_GBO0;
assign R14C3_GB00 = R14C4_GBO0;
assign R14C4_GB00 = R14C4_GBO0;
assign R14C5_GB00 = R14C4_GBO0;
assign R14C6_GB00 = R14C4_GBO0;
assign R15C2_GB00 = R15C4_GBO0;
assign R15C3_GB00 = R15C4_GBO0;
assign R15C4_GB00 = R15C4_GBO0;
assign R15C5_GB00 = R15C4_GBO0;
assign R15C6_GB00 = R15C4_GBO0;
assign R16C2_GB00 = R16C4_GBO0;
assign R16C3_GB00 = R16C4_GBO0;
assign R16C4_GB00 = R16C4_GBO0;
assign R16C5_GB00 = R16C4_GBO0;
assign R16C6_GB00 = R16C4_GBO0;
assign R17C2_GB00 = R17C4_GBO0;
assign R17C3_GB00 = R17C4_GBO0;
assign R17C4_GB00 = R17C4_GBO0;
assign R17C5_GB00 = R17C4_GBO0;
assign R17C6_GB00 = R17C4_GBO0;
assign R18C2_GB00 = R18C4_GBO0;
assign R18C3_GB00 = R18C4_GBO0;
assign R18C4_GB00 = R18C4_GBO0;
assign R18C5_GB00 = R18C4_GBO0;
assign R18C6_GB00 = R18C4_GBO0;
assign R20C2_GB00 = R20C4_GBO0;
assign R20C3_GB00 = R20C4_GBO0;
assign R20C4_GB00 = R20C4_GBO0;
assign R20C5_GB00 = R20C4_GBO0;
assign R20C6_GB00 = R20C4_GBO0;
assign R21C2_GB00 = R21C4_GBO0;
assign R21C3_GB00 = R21C4_GBO0;
assign R21C4_GB00 = R21C4_GBO0;
assign R21C5_GB00 = R21C4_GBO0;
assign R21C6_GB00 = R21C4_GBO0;
assign R22C2_GB00 = R22C4_GBO0;
assign R22C3_GB00 = R22C4_GBO0;
assign R22C4_GB00 = R22C4_GBO0;
assign R22C5_GB00 = R22C4_GBO0;
assign R22C6_GB00 = R22C4_GBO0;
assign R23C2_GB00 = R23C4_GBO0;
assign R23C3_GB00 = R23C4_GBO0;
assign R23C4_GB00 = R23C4_GBO0;
assign R23C5_GB00 = R23C4_GBO0;
assign R23C6_GB00 = R23C4_GBO0;
assign R24C2_GB00 = R24C4_GBO0;
assign R24C3_GB00 = R24C4_GBO0;
assign R24C4_GB00 = R24C4_GBO0;
assign R24C5_GB00 = R24C4_GBO0;
assign R24C6_GB00 = R24C4_GBO0;
assign R25C2_GB00 = R25C4_GBO0;
assign R25C3_GB00 = R25C4_GBO0;
assign R25C4_GB00 = R25C4_GBO0;
assign R25C5_GB00 = R25C4_GBO0;
assign R25C6_GB00 = R25C4_GBO0;
assign R26C2_GB00 = R26C4_GBO0;
assign R26C3_GB00 = R26C4_GBO0;
assign R26C4_GB00 = R26C4_GBO0;
assign R26C5_GB00 = R26C4_GBO0;
assign R26C6_GB00 = R26C4_GBO0;
assign R27C2_GB00 = R27C4_GBO0;
assign R27C3_GB00 = R27C4_GBO0;
assign R27C4_GB00 = R27C4_GBO0;
assign R27C5_GB00 = R27C4_GBO0;
assign R27C6_GB00 = R27C4_GBO0;
assign R11C9_GB00 = R11C8_GBO0;
assign R11C10_GB00 = R11C8_GBO0;
assign R11C7_GB00 = R11C8_GBO0;
assign R11C8_GB00 = R11C8_GBO0;
assign R12C9_GB00 = R12C8_GBO0;
assign R12C10_GB00 = R12C8_GBO0;
assign R12C7_GB00 = R12C8_GBO0;
assign R12C8_GB00 = R12C8_GBO0;
assign R13C9_GB00 = R13C8_GBO0;
assign R13C10_GB00 = R13C8_GBO0;
assign R13C7_GB00 = R13C8_GBO0;
assign R13C8_GB00 = R13C8_GBO0;
assign R14C9_GB00 = R14C8_GBO0;
assign R14C10_GB00 = R14C8_GBO0;
assign R14C7_GB00 = R14C8_GBO0;
assign R14C8_GB00 = R14C8_GBO0;
assign R15C9_GB00 = R15C8_GBO0;
assign R15C10_GB00 = R15C8_GBO0;
assign R15C7_GB00 = R15C8_GBO0;
assign R15C8_GB00 = R15C8_GBO0;
assign R16C9_GB00 = R16C8_GBO0;
assign R16C10_GB00 = R16C8_GBO0;
assign R16C7_GB00 = R16C8_GBO0;
assign R16C8_GB00 = R16C8_GBO0;
assign R17C9_GB00 = R17C8_GBO0;
assign R17C10_GB00 = R17C8_GBO0;
assign R17C7_GB00 = R17C8_GBO0;
assign R17C8_GB00 = R17C8_GBO0;
assign R18C9_GB00 = R18C8_GBO0;
assign R18C10_GB00 = R18C8_GBO0;
assign R18C7_GB00 = R18C8_GBO0;
assign R18C8_GB00 = R18C8_GBO0;
assign R20C9_GB00 = R20C8_GBO0;
assign R20C10_GB00 = R20C8_GBO0;
assign R20C7_GB00 = R20C8_GBO0;
assign R20C8_GB00 = R20C8_GBO0;
assign R21C9_GB00 = R21C8_GBO0;
assign R21C10_GB00 = R21C8_GBO0;
assign R21C7_GB00 = R21C8_GBO0;
assign R21C8_GB00 = R21C8_GBO0;
assign R22C9_GB00 = R22C8_GBO0;
assign R22C10_GB00 = R22C8_GBO0;
assign R22C7_GB00 = R22C8_GBO0;
assign R22C8_GB00 = R22C8_GBO0;
assign R23C9_GB00 = R23C8_GBO0;
assign R23C10_GB00 = R23C8_GBO0;
assign R23C7_GB00 = R23C8_GBO0;
assign R23C8_GB00 = R23C8_GBO0;
assign R24C9_GB00 = R24C8_GBO0;
assign R24C10_GB00 = R24C8_GBO0;
assign R24C7_GB00 = R24C8_GBO0;
assign R24C8_GB00 = R24C8_GBO0;
assign R25C9_GB00 = R25C8_GBO0;
assign R25C10_GB00 = R25C8_GBO0;
assign R25C7_GB00 = R25C8_GBO0;
assign R25C8_GB00 = R25C8_GBO0;
assign R26C9_GB00 = R26C8_GBO0;
assign R26C10_GB00 = R26C8_GBO0;
assign R26C7_GB00 = R26C8_GBO0;
assign R26C8_GB00 = R26C8_GBO0;
assign R27C9_GB00 = R27C8_GBO0;
assign R27C10_GB00 = R27C8_GBO0;
assign R27C7_GB00 = R27C8_GBO0;
assign R27C8_GB00 = R27C8_GBO0;
assign R11C11_GB00 = R11C12_GBO0;
assign R11C12_GB00 = R11C12_GBO0;
assign R11C13_GB00 = R11C12_GBO0;
assign R11C14_GB00 = R11C12_GBO0;
assign R12C11_GB00 = R12C12_GBO0;
assign R12C12_GB00 = R12C12_GBO0;
assign R12C13_GB00 = R12C12_GBO0;
assign R12C14_GB00 = R12C12_GBO0;
assign R13C11_GB00 = R13C12_GBO0;
assign R13C12_GB00 = R13C12_GBO0;
assign R13C13_GB00 = R13C12_GBO0;
assign R13C14_GB00 = R13C12_GBO0;
assign R14C11_GB00 = R14C12_GBO0;
assign R14C12_GB00 = R14C12_GBO0;
assign R14C13_GB00 = R14C12_GBO0;
assign R14C14_GB00 = R14C12_GBO0;
assign R15C11_GB00 = R15C12_GBO0;
assign R15C12_GB00 = R15C12_GBO0;
assign R15C13_GB00 = R15C12_GBO0;
assign R15C14_GB00 = R15C12_GBO0;
assign R16C11_GB00 = R16C12_GBO0;
assign R16C12_GB00 = R16C12_GBO0;
assign R16C13_GB00 = R16C12_GBO0;
assign R16C14_GB00 = R16C12_GBO0;
assign R17C11_GB00 = R17C12_GBO0;
assign R17C12_GB00 = R17C12_GBO0;
assign R17C13_GB00 = R17C12_GBO0;
assign R17C14_GB00 = R17C12_GBO0;
assign R18C11_GB00 = R18C12_GBO0;
assign R18C12_GB00 = R18C12_GBO0;
assign R18C13_GB00 = R18C12_GBO0;
assign R18C14_GB00 = R18C12_GBO0;
assign R20C11_GB00 = R20C12_GBO0;
assign R20C12_GB00 = R20C12_GBO0;
assign R20C13_GB00 = R20C12_GBO0;
assign R20C14_GB00 = R20C12_GBO0;
assign R21C11_GB00 = R21C12_GBO0;
assign R21C12_GB00 = R21C12_GBO0;
assign R21C13_GB00 = R21C12_GBO0;
assign R21C14_GB00 = R21C12_GBO0;
assign R22C11_GB00 = R22C12_GBO0;
assign R22C12_GB00 = R22C12_GBO0;
assign R22C13_GB00 = R22C12_GBO0;
assign R22C14_GB00 = R22C12_GBO0;
assign R23C11_GB00 = R23C12_GBO0;
assign R23C12_GB00 = R23C12_GBO0;
assign R23C13_GB00 = R23C12_GBO0;
assign R23C14_GB00 = R23C12_GBO0;
assign R24C11_GB00 = R24C12_GBO0;
assign R24C12_GB00 = R24C12_GBO0;
assign R24C13_GB00 = R24C12_GBO0;
assign R24C14_GB00 = R24C12_GBO0;
assign R25C11_GB00 = R25C12_GBO0;
assign R25C12_GB00 = R25C12_GBO0;
assign R25C13_GB00 = R25C12_GBO0;
assign R25C14_GB00 = R25C12_GBO0;
assign R26C11_GB00 = R26C12_GBO0;
assign R26C12_GB00 = R26C12_GBO0;
assign R26C13_GB00 = R26C12_GBO0;
assign R26C14_GB00 = R26C12_GBO0;
assign R27C11_GB00 = R27C12_GBO0;
assign R27C12_GB00 = R27C12_GBO0;
assign R27C13_GB00 = R27C12_GBO0;
assign R27C14_GB00 = R27C12_GBO0;
assign R11C17_GB00 = R11C16_GBO0;
assign R11C18_GB00 = R11C16_GBO0;
assign R11C15_GB00 = R11C16_GBO0;
assign R11C16_GB00 = R11C16_GBO0;
assign R12C17_GB00 = R12C16_GBO0;
assign R12C18_GB00 = R12C16_GBO0;
assign R12C15_GB00 = R12C16_GBO0;
assign R12C16_GB00 = R12C16_GBO0;
assign R13C17_GB00 = R13C16_GBO0;
assign R13C18_GB00 = R13C16_GBO0;
assign R13C15_GB00 = R13C16_GBO0;
assign R13C16_GB00 = R13C16_GBO0;
assign R14C17_GB00 = R14C16_GBO0;
assign R14C18_GB00 = R14C16_GBO0;
assign R14C15_GB00 = R14C16_GBO0;
assign R14C16_GB00 = R14C16_GBO0;
assign R15C17_GB00 = R15C16_GBO0;
assign R15C18_GB00 = R15C16_GBO0;
assign R15C15_GB00 = R15C16_GBO0;
assign R15C16_GB00 = R15C16_GBO0;
assign R16C17_GB00 = R16C16_GBO0;
assign R16C18_GB00 = R16C16_GBO0;
assign R16C15_GB00 = R16C16_GBO0;
assign R16C16_GB00 = R16C16_GBO0;
assign R17C17_GB00 = R17C16_GBO0;
assign R17C18_GB00 = R17C16_GBO0;
assign R17C15_GB00 = R17C16_GBO0;
assign R17C16_GB00 = R17C16_GBO0;
assign R18C17_GB00 = R18C16_GBO0;
assign R18C18_GB00 = R18C16_GBO0;
assign R18C15_GB00 = R18C16_GBO0;
assign R18C16_GB00 = R18C16_GBO0;
assign R20C17_GB00 = R20C16_GBO0;
assign R20C18_GB00 = R20C16_GBO0;
assign R20C15_GB00 = R20C16_GBO0;
assign R20C16_GB00 = R20C16_GBO0;
assign R21C17_GB00 = R21C16_GBO0;
assign R21C18_GB00 = R21C16_GBO0;
assign R21C15_GB00 = R21C16_GBO0;
assign R21C16_GB00 = R21C16_GBO0;
assign R22C17_GB00 = R22C16_GBO0;
assign R22C18_GB00 = R22C16_GBO0;
assign R22C15_GB00 = R22C16_GBO0;
assign R22C16_GB00 = R22C16_GBO0;
assign R23C17_GB00 = R23C16_GBO0;
assign R23C18_GB00 = R23C16_GBO0;
assign R23C15_GB00 = R23C16_GBO0;
assign R23C16_GB00 = R23C16_GBO0;
assign R24C17_GB00 = R24C16_GBO0;
assign R24C18_GB00 = R24C16_GBO0;
assign R24C15_GB00 = R24C16_GBO0;
assign R24C16_GB00 = R24C16_GBO0;
assign R25C17_GB00 = R25C16_GBO0;
assign R25C18_GB00 = R25C16_GBO0;
assign R25C15_GB00 = R25C16_GBO0;
assign R25C16_GB00 = R25C16_GBO0;
assign R26C17_GB00 = R26C16_GBO0;
assign R26C18_GB00 = R26C16_GBO0;
assign R26C15_GB00 = R26C16_GBO0;
assign R26C16_GB00 = R26C16_GBO0;
assign R27C17_GB00 = R27C16_GBO0;
assign R27C18_GB00 = R27C16_GBO0;
assign R27C15_GB00 = R27C16_GBO0;
assign R27C16_GB00 = R27C16_GBO0;
assign R11C19_GB00 = R11C20_GBO0;
assign R11C20_GB00 = R11C20_GBO0;
assign R11C21_GB00 = R11C20_GBO0;
assign R11C22_GB00 = R11C20_GBO0;
assign R12C19_GB00 = R12C20_GBO0;
assign R12C20_GB00 = R12C20_GBO0;
assign R12C21_GB00 = R12C20_GBO0;
assign R12C22_GB00 = R12C20_GBO0;
assign R13C19_GB00 = R13C20_GBO0;
assign R13C20_GB00 = R13C20_GBO0;
assign R13C21_GB00 = R13C20_GBO0;
assign R13C22_GB00 = R13C20_GBO0;
assign R14C19_GB00 = R14C20_GBO0;
assign R14C20_GB00 = R14C20_GBO0;
assign R14C21_GB00 = R14C20_GBO0;
assign R14C22_GB00 = R14C20_GBO0;
assign R15C19_GB00 = R15C20_GBO0;
assign R15C20_GB00 = R15C20_GBO0;
assign R15C21_GB00 = R15C20_GBO0;
assign R15C22_GB00 = R15C20_GBO0;
assign R16C19_GB00 = R16C20_GBO0;
assign R16C20_GB00 = R16C20_GBO0;
assign R16C21_GB00 = R16C20_GBO0;
assign R16C22_GB00 = R16C20_GBO0;
assign R17C19_GB00 = R17C20_GBO0;
assign R17C20_GB00 = R17C20_GBO0;
assign R17C21_GB00 = R17C20_GBO0;
assign R17C22_GB00 = R17C20_GBO0;
assign R18C19_GB00 = R18C20_GBO0;
assign R18C20_GB00 = R18C20_GBO0;
assign R18C21_GB00 = R18C20_GBO0;
assign R18C22_GB00 = R18C20_GBO0;
assign R20C19_GB00 = R20C20_GBO0;
assign R20C20_GB00 = R20C20_GBO0;
assign R20C21_GB00 = R20C20_GBO0;
assign R20C22_GB00 = R20C20_GBO0;
assign R21C19_GB00 = R21C20_GBO0;
assign R21C20_GB00 = R21C20_GBO0;
assign R21C21_GB00 = R21C20_GBO0;
assign R21C22_GB00 = R21C20_GBO0;
assign R22C19_GB00 = R22C20_GBO0;
assign R22C20_GB00 = R22C20_GBO0;
assign R22C21_GB00 = R22C20_GBO0;
assign R22C22_GB00 = R22C20_GBO0;
assign R23C19_GB00 = R23C20_GBO0;
assign R23C20_GB00 = R23C20_GBO0;
assign R23C21_GB00 = R23C20_GBO0;
assign R23C22_GB00 = R23C20_GBO0;
assign R24C19_GB00 = R24C20_GBO0;
assign R24C20_GB00 = R24C20_GBO0;
assign R24C21_GB00 = R24C20_GBO0;
assign R24C22_GB00 = R24C20_GBO0;
assign R25C19_GB00 = R25C20_GBO0;
assign R25C20_GB00 = R25C20_GBO0;
assign R25C21_GB00 = R25C20_GBO0;
assign R25C22_GB00 = R25C20_GBO0;
assign R26C19_GB00 = R26C20_GBO0;
assign R26C20_GB00 = R26C20_GBO0;
assign R26C21_GB00 = R26C20_GBO0;
assign R26C22_GB00 = R26C20_GBO0;
assign R27C19_GB00 = R27C20_GBO0;
assign R27C20_GB00 = R27C20_GBO0;
assign R27C21_GB00 = R27C20_GBO0;
assign R27C22_GB00 = R27C20_GBO0;
assign R11C23_GB00 = R11C24_GBO0;
assign R11C24_GB00 = R11C24_GBO0;
assign R11C25_GB00 = R11C24_GBO0;
assign R11C26_GB00 = R11C24_GBO0;
assign R11C27_GB00 = R11C24_GBO0;
assign R11C28_GB00 = R11C24_GBO0;
assign R12C23_GB00 = R12C24_GBO0;
assign R12C24_GB00 = R12C24_GBO0;
assign R12C25_GB00 = R12C24_GBO0;
assign R12C26_GB00 = R12C24_GBO0;
assign R12C27_GB00 = R12C24_GBO0;
assign R12C28_GB00 = R12C24_GBO0;
assign R13C23_GB00 = R13C24_GBO0;
assign R13C24_GB00 = R13C24_GBO0;
assign R13C25_GB00 = R13C24_GBO0;
assign R13C26_GB00 = R13C24_GBO0;
assign R13C27_GB00 = R13C24_GBO0;
assign R13C28_GB00 = R13C24_GBO0;
assign R14C23_GB00 = R14C24_GBO0;
assign R14C24_GB00 = R14C24_GBO0;
assign R14C25_GB00 = R14C24_GBO0;
assign R14C26_GB00 = R14C24_GBO0;
assign R14C27_GB00 = R14C24_GBO0;
assign R14C28_GB00 = R14C24_GBO0;
assign R15C23_GB00 = R15C24_GBO0;
assign R15C24_GB00 = R15C24_GBO0;
assign R15C25_GB00 = R15C24_GBO0;
assign R15C26_GB00 = R15C24_GBO0;
assign R15C27_GB00 = R15C24_GBO0;
assign R15C28_GB00 = R15C24_GBO0;
assign R16C23_GB00 = R16C24_GBO0;
assign R16C24_GB00 = R16C24_GBO0;
assign R16C25_GB00 = R16C24_GBO0;
assign R16C26_GB00 = R16C24_GBO0;
assign R16C27_GB00 = R16C24_GBO0;
assign R16C28_GB00 = R16C24_GBO0;
assign R17C23_GB00 = R17C24_GBO0;
assign R17C24_GB00 = R17C24_GBO0;
assign R17C25_GB00 = R17C24_GBO0;
assign R17C26_GB00 = R17C24_GBO0;
assign R17C27_GB00 = R17C24_GBO0;
assign R17C28_GB00 = R17C24_GBO0;
assign R18C23_GB00 = R18C24_GBO0;
assign R18C24_GB00 = R18C24_GBO0;
assign R18C25_GB00 = R18C24_GBO0;
assign R18C26_GB00 = R18C24_GBO0;
assign R18C27_GB00 = R18C24_GBO0;
assign R18C28_GB00 = R18C24_GBO0;
assign R20C23_GB00 = R20C24_GBO0;
assign R20C24_GB00 = R20C24_GBO0;
assign R20C25_GB00 = R20C24_GBO0;
assign R20C26_GB00 = R20C24_GBO0;
assign R20C27_GB00 = R20C24_GBO0;
assign R20C28_GB00 = R20C24_GBO0;
assign R21C23_GB00 = R21C24_GBO0;
assign R21C24_GB00 = R21C24_GBO0;
assign R21C25_GB00 = R21C24_GBO0;
assign R21C26_GB00 = R21C24_GBO0;
assign R21C27_GB00 = R21C24_GBO0;
assign R21C28_GB00 = R21C24_GBO0;
assign R22C23_GB00 = R22C24_GBO0;
assign R22C24_GB00 = R22C24_GBO0;
assign R22C25_GB00 = R22C24_GBO0;
assign R22C26_GB00 = R22C24_GBO0;
assign R22C27_GB00 = R22C24_GBO0;
assign R22C28_GB00 = R22C24_GBO0;
assign R23C23_GB00 = R23C24_GBO0;
assign R23C24_GB00 = R23C24_GBO0;
assign R23C25_GB00 = R23C24_GBO0;
assign R23C26_GB00 = R23C24_GBO0;
assign R23C27_GB00 = R23C24_GBO0;
assign R23C28_GB00 = R23C24_GBO0;
assign R24C23_GB00 = R24C24_GBO0;
assign R24C24_GB00 = R24C24_GBO0;
assign R24C25_GB00 = R24C24_GBO0;
assign R24C26_GB00 = R24C24_GBO0;
assign R24C27_GB00 = R24C24_GBO0;
assign R24C28_GB00 = R24C24_GBO0;
assign R25C23_GB00 = R25C24_GBO0;
assign R25C24_GB00 = R25C24_GBO0;
assign R25C25_GB00 = R25C24_GBO0;
assign R25C26_GB00 = R25C24_GBO0;
assign R25C27_GB00 = R25C24_GBO0;
assign R25C28_GB00 = R25C24_GBO0;
assign R26C23_GB00 = R26C24_GBO0;
assign R26C24_GB00 = R26C24_GBO0;
assign R26C25_GB00 = R26C24_GBO0;
assign R26C26_GB00 = R26C24_GBO0;
assign R26C27_GB00 = R26C24_GBO0;
assign R26C28_GB00 = R26C24_GBO0;
assign R27C23_GB00 = R27C24_GBO0;
assign R27C24_GB00 = R27C24_GBO0;
assign R27C25_GB00 = R27C24_GBO0;
assign R27C26_GB00 = R27C24_GBO0;
assign R27C27_GB00 = R27C24_GBO0;
assign R27C28_GB00 = R27C24_GBO0;
assign R11C2_GB10 = R11C3_GBO0;
assign R11C3_GB10 = R11C3_GBO0;
assign R11C4_GB10 = R11C3_GBO0;
assign R11C5_GB10 = R11C3_GBO0;
assign R12C2_GB10 = R12C3_GBO0;
assign R12C3_GB10 = R12C3_GBO0;
assign R12C4_GB10 = R12C3_GBO0;
assign R12C5_GB10 = R12C3_GBO0;
assign R13C2_GB10 = R13C3_GBO0;
assign R13C3_GB10 = R13C3_GBO0;
assign R13C4_GB10 = R13C3_GBO0;
assign R13C5_GB10 = R13C3_GBO0;
assign R14C2_GB10 = R14C3_GBO0;
assign R14C3_GB10 = R14C3_GBO0;
assign R14C4_GB10 = R14C3_GBO0;
assign R14C5_GB10 = R14C3_GBO0;
assign R15C2_GB10 = R15C3_GBO0;
assign R15C3_GB10 = R15C3_GBO0;
assign R15C4_GB10 = R15C3_GBO0;
assign R15C5_GB10 = R15C3_GBO0;
assign R16C2_GB10 = R16C3_GBO0;
assign R16C3_GB10 = R16C3_GBO0;
assign R16C4_GB10 = R16C3_GBO0;
assign R16C5_GB10 = R16C3_GBO0;
assign R17C2_GB10 = R17C3_GBO0;
assign R17C3_GB10 = R17C3_GBO0;
assign R17C4_GB10 = R17C3_GBO0;
assign R17C5_GB10 = R17C3_GBO0;
assign R18C2_GB10 = R18C3_GBO0;
assign R18C3_GB10 = R18C3_GBO0;
assign R18C4_GB10 = R18C3_GBO0;
assign R18C5_GB10 = R18C3_GBO0;
assign R20C2_GB10 = R20C3_GBO0;
assign R20C3_GB10 = R20C3_GBO0;
assign R20C4_GB10 = R20C3_GBO0;
assign R20C5_GB10 = R20C3_GBO0;
assign R21C2_GB10 = R21C3_GBO0;
assign R21C3_GB10 = R21C3_GBO0;
assign R21C4_GB10 = R21C3_GBO0;
assign R21C5_GB10 = R21C3_GBO0;
assign R22C2_GB10 = R22C3_GBO0;
assign R22C3_GB10 = R22C3_GBO0;
assign R22C4_GB10 = R22C3_GBO0;
assign R22C5_GB10 = R22C3_GBO0;
assign R23C2_GB10 = R23C3_GBO0;
assign R23C3_GB10 = R23C3_GBO0;
assign R23C4_GB10 = R23C3_GBO0;
assign R23C5_GB10 = R23C3_GBO0;
assign R24C2_GB10 = R24C3_GBO0;
assign R24C3_GB10 = R24C3_GBO0;
assign R24C4_GB10 = R24C3_GBO0;
assign R24C5_GB10 = R24C3_GBO0;
assign R25C2_GB10 = R25C3_GBO0;
assign R25C3_GB10 = R25C3_GBO0;
assign R25C4_GB10 = R25C3_GBO0;
assign R25C5_GB10 = R25C3_GBO0;
assign R26C2_GB10 = R26C3_GBO0;
assign R26C3_GB10 = R26C3_GBO0;
assign R26C4_GB10 = R26C3_GBO0;
assign R26C5_GB10 = R26C3_GBO0;
assign R27C2_GB10 = R27C3_GBO0;
assign R27C3_GB10 = R27C3_GBO0;
assign R27C4_GB10 = R27C3_GBO0;
assign R27C5_GB10 = R27C3_GBO0;
assign R11C9_GB10 = R11C7_GBO0;
assign R11C6_GB10 = R11C7_GBO0;
assign R11C7_GB10 = R11C7_GBO0;
assign R11C8_GB10 = R11C7_GBO0;
assign R12C9_GB10 = R12C7_GBO0;
assign R12C6_GB10 = R12C7_GBO0;
assign R12C7_GB10 = R12C7_GBO0;
assign R12C8_GB10 = R12C7_GBO0;
assign R13C9_GB10 = R13C7_GBO0;
assign R13C6_GB10 = R13C7_GBO0;
assign R13C7_GB10 = R13C7_GBO0;
assign R13C8_GB10 = R13C7_GBO0;
assign R14C9_GB10 = R14C7_GBO0;
assign R14C6_GB10 = R14C7_GBO0;
assign R14C7_GB10 = R14C7_GBO0;
assign R14C8_GB10 = R14C7_GBO0;
assign R15C9_GB10 = R15C7_GBO0;
assign R15C6_GB10 = R15C7_GBO0;
assign R15C7_GB10 = R15C7_GBO0;
assign R15C8_GB10 = R15C7_GBO0;
assign R16C9_GB10 = R16C7_GBO0;
assign R16C6_GB10 = R16C7_GBO0;
assign R16C7_GB10 = R16C7_GBO0;
assign R16C8_GB10 = R16C7_GBO0;
assign R17C9_GB10 = R17C7_GBO0;
assign R17C6_GB10 = R17C7_GBO0;
assign R17C7_GB10 = R17C7_GBO0;
assign R17C8_GB10 = R17C7_GBO0;
assign R18C9_GB10 = R18C7_GBO0;
assign R18C6_GB10 = R18C7_GBO0;
assign R18C7_GB10 = R18C7_GBO0;
assign R18C8_GB10 = R18C7_GBO0;
assign R20C9_GB10 = R20C7_GBO0;
assign R20C6_GB10 = R20C7_GBO0;
assign R20C7_GB10 = R20C7_GBO0;
assign R20C8_GB10 = R20C7_GBO0;
assign R21C9_GB10 = R21C7_GBO0;
assign R21C6_GB10 = R21C7_GBO0;
assign R21C7_GB10 = R21C7_GBO0;
assign R21C8_GB10 = R21C7_GBO0;
assign R22C9_GB10 = R22C7_GBO0;
assign R22C6_GB10 = R22C7_GBO0;
assign R22C7_GB10 = R22C7_GBO0;
assign R22C8_GB10 = R22C7_GBO0;
assign R23C9_GB10 = R23C7_GBO0;
assign R23C6_GB10 = R23C7_GBO0;
assign R23C7_GB10 = R23C7_GBO0;
assign R23C8_GB10 = R23C7_GBO0;
assign R24C9_GB10 = R24C7_GBO0;
assign R24C6_GB10 = R24C7_GBO0;
assign R24C7_GB10 = R24C7_GBO0;
assign R24C8_GB10 = R24C7_GBO0;
assign R25C9_GB10 = R25C7_GBO0;
assign R25C6_GB10 = R25C7_GBO0;
assign R25C7_GB10 = R25C7_GBO0;
assign R25C8_GB10 = R25C7_GBO0;
assign R26C9_GB10 = R26C7_GBO0;
assign R26C6_GB10 = R26C7_GBO0;
assign R26C7_GB10 = R26C7_GBO0;
assign R26C8_GB10 = R26C7_GBO0;
assign R27C9_GB10 = R27C7_GBO0;
assign R27C6_GB10 = R27C7_GBO0;
assign R27C7_GB10 = R27C7_GBO0;
assign R27C8_GB10 = R27C7_GBO0;
assign R11C10_GB10 = R11C11_GBO0;
assign R11C11_GB10 = R11C11_GBO0;
assign R11C12_GB10 = R11C11_GBO0;
assign R11C13_GB10 = R11C11_GBO0;
assign R12C10_GB10 = R12C11_GBO0;
assign R12C11_GB10 = R12C11_GBO0;
assign R12C12_GB10 = R12C11_GBO0;
assign R12C13_GB10 = R12C11_GBO0;
assign R13C10_GB10 = R13C11_GBO0;
assign R13C11_GB10 = R13C11_GBO0;
assign R13C12_GB10 = R13C11_GBO0;
assign R13C13_GB10 = R13C11_GBO0;
assign R14C10_GB10 = R14C11_GBO0;
assign R14C11_GB10 = R14C11_GBO0;
assign R14C12_GB10 = R14C11_GBO0;
assign R14C13_GB10 = R14C11_GBO0;
assign R15C10_GB10 = R15C11_GBO0;
assign R15C11_GB10 = R15C11_GBO0;
assign R15C12_GB10 = R15C11_GBO0;
assign R15C13_GB10 = R15C11_GBO0;
assign R16C10_GB10 = R16C11_GBO0;
assign R16C11_GB10 = R16C11_GBO0;
assign R16C12_GB10 = R16C11_GBO0;
assign R16C13_GB10 = R16C11_GBO0;
assign R17C10_GB10 = R17C11_GBO0;
assign R17C11_GB10 = R17C11_GBO0;
assign R17C12_GB10 = R17C11_GBO0;
assign R17C13_GB10 = R17C11_GBO0;
assign R18C10_GB10 = R18C11_GBO0;
assign R18C11_GB10 = R18C11_GBO0;
assign R18C12_GB10 = R18C11_GBO0;
assign R18C13_GB10 = R18C11_GBO0;
assign R20C10_GB10 = R20C11_GBO0;
assign R20C11_GB10 = R20C11_GBO0;
assign R20C12_GB10 = R20C11_GBO0;
assign R20C13_GB10 = R20C11_GBO0;
assign R21C10_GB10 = R21C11_GBO0;
assign R21C11_GB10 = R21C11_GBO0;
assign R21C12_GB10 = R21C11_GBO0;
assign R21C13_GB10 = R21C11_GBO0;
assign R22C10_GB10 = R22C11_GBO0;
assign R22C11_GB10 = R22C11_GBO0;
assign R22C12_GB10 = R22C11_GBO0;
assign R22C13_GB10 = R22C11_GBO0;
assign R23C10_GB10 = R23C11_GBO0;
assign R23C11_GB10 = R23C11_GBO0;
assign R23C12_GB10 = R23C11_GBO0;
assign R23C13_GB10 = R23C11_GBO0;
assign R24C10_GB10 = R24C11_GBO0;
assign R24C11_GB10 = R24C11_GBO0;
assign R24C12_GB10 = R24C11_GBO0;
assign R24C13_GB10 = R24C11_GBO0;
assign R25C10_GB10 = R25C11_GBO0;
assign R25C11_GB10 = R25C11_GBO0;
assign R25C12_GB10 = R25C11_GBO0;
assign R25C13_GB10 = R25C11_GBO0;
assign R26C10_GB10 = R26C11_GBO0;
assign R26C11_GB10 = R26C11_GBO0;
assign R26C12_GB10 = R26C11_GBO0;
assign R26C13_GB10 = R26C11_GBO0;
assign R27C10_GB10 = R27C11_GBO0;
assign R27C11_GB10 = R27C11_GBO0;
assign R27C12_GB10 = R27C11_GBO0;
assign R27C13_GB10 = R27C11_GBO0;
assign R11C17_GB10 = R11C15_GBO0;
assign R11C14_GB10 = R11C15_GBO0;
assign R11C15_GB10 = R11C15_GBO0;
assign R11C16_GB10 = R11C15_GBO0;
assign R12C17_GB10 = R12C15_GBO0;
assign R12C14_GB10 = R12C15_GBO0;
assign R12C15_GB10 = R12C15_GBO0;
assign R12C16_GB10 = R12C15_GBO0;
assign R13C17_GB10 = R13C15_GBO0;
assign R13C14_GB10 = R13C15_GBO0;
assign R13C15_GB10 = R13C15_GBO0;
assign R13C16_GB10 = R13C15_GBO0;
assign R14C17_GB10 = R14C15_GBO0;
assign R14C14_GB10 = R14C15_GBO0;
assign R14C15_GB10 = R14C15_GBO0;
assign R14C16_GB10 = R14C15_GBO0;
assign R15C17_GB10 = R15C15_GBO0;
assign R15C14_GB10 = R15C15_GBO0;
assign R15C15_GB10 = R15C15_GBO0;
assign R15C16_GB10 = R15C15_GBO0;
assign R16C17_GB10 = R16C15_GBO0;
assign R16C14_GB10 = R16C15_GBO0;
assign R16C15_GB10 = R16C15_GBO0;
assign R16C16_GB10 = R16C15_GBO0;
assign R17C17_GB10 = R17C15_GBO0;
assign R17C14_GB10 = R17C15_GBO0;
assign R17C15_GB10 = R17C15_GBO0;
assign R17C16_GB10 = R17C15_GBO0;
assign R18C17_GB10 = R18C15_GBO0;
assign R18C14_GB10 = R18C15_GBO0;
assign R18C15_GB10 = R18C15_GBO0;
assign R18C16_GB10 = R18C15_GBO0;
assign R20C17_GB10 = R20C15_GBO0;
assign R20C14_GB10 = R20C15_GBO0;
assign R20C15_GB10 = R20C15_GBO0;
assign R20C16_GB10 = R20C15_GBO0;
assign R21C17_GB10 = R21C15_GBO0;
assign R21C14_GB10 = R21C15_GBO0;
assign R21C15_GB10 = R21C15_GBO0;
assign R21C16_GB10 = R21C15_GBO0;
assign R22C17_GB10 = R22C15_GBO0;
assign R22C14_GB10 = R22C15_GBO0;
assign R22C15_GB10 = R22C15_GBO0;
assign R22C16_GB10 = R22C15_GBO0;
assign R23C17_GB10 = R23C15_GBO0;
assign R23C14_GB10 = R23C15_GBO0;
assign R23C15_GB10 = R23C15_GBO0;
assign R23C16_GB10 = R23C15_GBO0;
assign R24C17_GB10 = R24C15_GBO0;
assign R24C14_GB10 = R24C15_GBO0;
assign R24C15_GB10 = R24C15_GBO0;
assign R24C16_GB10 = R24C15_GBO0;
assign R25C17_GB10 = R25C15_GBO0;
assign R25C14_GB10 = R25C15_GBO0;
assign R25C15_GB10 = R25C15_GBO0;
assign R25C16_GB10 = R25C15_GBO0;
assign R26C17_GB10 = R26C15_GBO0;
assign R26C14_GB10 = R26C15_GBO0;
assign R26C15_GB10 = R26C15_GBO0;
assign R26C16_GB10 = R26C15_GBO0;
assign R27C17_GB10 = R27C15_GBO0;
assign R27C14_GB10 = R27C15_GBO0;
assign R27C15_GB10 = R27C15_GBO0;
assign R27C16_GB10 = R27C15_GBO0;
assign R11C18_GB10 = R11C19_GBO0;
assign R11C19_GB10 = R11C19_GBO0;
assign R11C20_GB10 = R11C19_GBO0;
assign R11C21_GB10 = R11C19_GBO0;
assign R12C18_GB10 = R12C19_GBO0;
assign R12C19_GB10 = R12C19_GBO0;
assign R12C20_GB10 = R12C19_GBO0;
assign R12C21_GB10 = R12C19_GBO0;
assign R13C18_GB10 = R13C19_GBO0;
assign R13C19_GB10 = R13C19_GBO0;
assign R13C20_GB10 = R13C19_GBO0;
assign R13C21_GB10 = R13C19_GBO0;
assign R14C18_GB10 = R14C19_GBO0;
assign R14C19_GB10 = R14C19_GBO0;
assign R14C20_GB10 = R14C19_GBO0;
assign R14C21_GB10 = R14C19_GBO0;
assign R15C18_GB10 = R15C19_GBO0;
assign R15C19_GB10 = R15C19_GBO0;
assign R15C20_GB10 = R15C19_GBO0;
assign R15C21_GB10 = R15C19_GBO0;
assign R16C18_GB10 = R16C19_GBO0;
assign R16C19_GB10 = R16C19_GBO0;
assign R16C20_GB10 = R16C19_GBO0;
assign R16C21_GB10 = R16C19_GBO0;
assign R17C18_GB10 = R17C19_GBO0;
assign R17C19_GB10 = R17C19_GBO0;
assign R17C20_GB10 = R17C19_GBO0;
assign R17C21_GB10 = R17C19_GBO0;
assign R18C18_GB10 = R18C19_GBO0;
assign R18C19_GB10 = R18C19_GBO0;
assign R18C20_GB10 = R18C19_GBO0;
assign R18C21_GB10 = R18C19_GBO0;
assign R20C18_GB10 = R20C19_GBO0;
assign R20C19_GB10 = R20C19_GBO0;
assign R20C20_GB10 = R20C19_GBO0;
assign R20C21_GB10 = R20C19_GBO0;
assign R21C18_GB10 = R21C19_GBO0;
assign R21C19_GB10 = R21C19_GBO0;
assign R21C20_GB10 = R21C19_GBO0;
assign R21C21_GB10 = R21C19_GBO0;
assign R22C18_GB10 = R22C19_GBO0;
assign R22C19_GB10 = R22C19_GBO0;
assign R22C20_GB10 = R22C19_GBO0;
assign R22C21_GB10 = R22C19_GBO0;
assign R23C18_GB10 = R23C19_GBO0;
assign R23C19_GB10 = R23C19_GBO0;
assign R23C20_GB10 = R23C19_GBO0;
assign R23C21_GB10 = R23C19_GBO0;
assign R24C18_GB10 = R24C19_GBO0;
assign R24C19_GB10 = R24C19_GBO0;
assign R24C20_GB10 = R24C19_GBO0;
assign R24C21_GB10 = R24C19_GBO0;
assign R25C18_GB10 = R25C19_GBO0;
assign R25C19_GB10 = R25C19_GBO0;
assign R25C20_GB10 = R25C19_GBO0;
assign R25C21_GB10 = R25C19_GBO0;
assign R26C18_GB10 = R26C19_GBO0;
assign R26C19_GB10 = R26C19_GBO0;
assign R26C20_GB10 = R26C19_GBO0;
assign R26C21_GB10 = R26C19_GBO0;
assign R27C18_GB10 = R27C19_GBO0;
assign R27C19_GB10 = R27C19_GBO0;
assign R27C20_GB10 = R27C19_GBO0;
assign R27C21_GB10 = R27C19_GBO0;
assign R11C25_GB10 = R11C23_GBO0;
assign R11C22_GB10 = R11C23_GBO0;
assign R11C23_GB10 = R11C23_GBO0;
assign R11C24_GB10 = R11C23_GBO0;
assign R12C25_GB10 = R12C23_GBO0;
assign R12C22_GB10 = R12C23_GBO0;
assign R12C23_GB10 = R12C23_GBO0;
assign R12C24_GB10 = R12C23_GBO0;
assign R13C25_GB10 = R13C23_GBO0;
assign R13C22_GB10 = R13C23_GBO0;
assign R13C23_GB10 = R13C23_GBO0;
assign R13C24_GB10 = R13C23_GBO0;
assign R14C25_GB10 = R14C23_GBO0;
assign R14C22_GB10 = R14C23_GBO0;
assign R14C23_GB10 = R14C23_GBO0;
assign R14C24_GB10 = R14C23_GBO0;
assign R15C25_GB10 = R15C23_GBO0;
assign R15C22_GB10 = R15C23_GBO0;
assign R15C23_GB10 = R15C23_GBO0;
assign R15C24_GB10 = R15C23_GBO0;
assign R16C25_GB10 = R16C23_GBO0;
assign R16C22_GB10 = R16C23_GBO0;
assign R16C23_GB10 = R16C23_GBO0;
assign R16C24_GB10 = R16C23_GBO0;
assign R17C25_GB10 = R17C23_GBO0;
assign R17C22_GB10 = R17C23_GBO0;
assign R17C23_GB10 = R17C23_GBO0;
assign R17C24_GB10 = R17C23_GBO0;
assign R18C25_GB10 = R18C23_GBO0;
assign R18C22_GB10 = R18C23_GBO0;
assign R18C23_GB10 = R18C23_GBO0;
assign R18C24_GB10 = R18C23_GBO0;
assign R20C25_GB10 = R20C23_GBO0;
assign R20C22_GB10 = R20C23_GBO0;
assign R20C23_GB10 = R20C23_GBO0;
assign R20C24_GB10 = R20C23_GBO0;
assign R21C25_GB10 = R21C23_GBO0;
assign R21C22_GB10 = R21C23_GBO0;
assign R21C23_GB10 = R21C23_GBO0;
assign R21C24_GB10 = R21C23_GBO0;
assign R22C25_GB10 = R22C23_GBO0;
assign R22C22_GB10 = R22C23_GBO0;
assign R22C23_GB10 = R22C23_GBO0;
assign R22C24_GB10 = R22C23_GBO0;
assign R23C25_GB10 = R23C23_GBO0;
assign R23C22_GB10 = R23C23_GBO0;
assign R23C23_GB10 = R23C23_GBO0;
assign R23C24_GB10 = R23C23_GBO0;
assign R24C25_GB10 = R24C23_GBO0;
assign R24C22_GB10 = R24C23_GBO0;
assign R24C23_GB10 = R24C23_GBO0;
assign R24C24_GB10 = R24C23_GBO0;
assign R25C25_GB10 = R25C23_GBO0;
assign R25C22_GB10 = R25C23_GBO0;
assign R25C23_GB10 = R25C23_GBO0;
assign R25C24_GB10 = R25C23_GBO0;
assign R26C25_GB10 = R26C23_GBO0;
assign R26C22_GB10 = R26C23_GBO0;
assign R26C23_GB10 = R26C23_GBO0;
assign R26C24_GB10 = R26C23_GBO0;
assign R27C25_GB10 = R27C23_GBO0;
assign R27C22_GB10 = R27C23_GBO0;
assign R27C23_GB10 = R27C23_GBO0;
assign R27C24_GB10 = R27C23_GBO0;
assign R11C26_GB10 = R11C27_GBO0;
assign R11C27_GB10 = R11C27_GBO0;
assign R11C28_GB10 = R11C27_GBO0;
assign R12C26_GB10 = R12C27_GBO0;
assign R12C27_GB10 = R12C27_GBO0;
assign R12C28_GB10 = R12C27_GBO0;
assign R13C26_GB10 = R13C27_GBO0;
assign R13C27_GB10 = R13C27_GBO0;
assign R13C28_GB10 = R13C27_GBO0;
assign R14C26_GB10 = R14C27_GBO0;
assign R14C27_GB10 = R14C27_GBO0;
assign R14C28_GB10 = R14C27_GBO0;
assign R15C26_GB10 = R15C27_GBO0;
assign R15C27_GB10 = R15C27_GBO0;
assign R15C28_GB10 = R15C27_GBO0;
assign R16C26_GB10 = R16C27_GBO0;
assign R16C27_GB10 = R16C27_GBO0;
assign R16C28_GB10 = R16C27_GBO0;
assign R17C26_GB10 = R17C27_GBO0;
assign R17C27_GB10 = R17C27_GBO0;
assign R17C28_GB10 = R17C27_GBO0;
assign R18C26_GB10 = R18C27_GBO0;
assign R18C27_GB10 = R18C27_GBO0;
assign R18C28_GB10 = R18C27_GBO0;
assign R20C26_GB10 = R20C27_GBO0;
assign R20C27_GB10 = R20C27_GBO0;
assign R20C28_GB10 = R20C27_GBO0;
assign R21C26_GB10 = R21C27_GBO0;
assign R21C27_GB10 = R21C27_GBO0;
assign R21C28_GB10 = R21C27_GBO0;
assign R22C26_GB10 = R22C27_GBO0;
assign R22C27_GB10 = R22C27_GBO0;
assign R22C28_GB10 = R22C27_GBO0;
assign R23C26_GB10 = R23C27_GBO0;
assign R23C27_GB10 = R23C27_GBO0;
assign R23C28_GB10 = R23C27_GBO0;
assign R24C26_GB10 = R24C27_GBO0;
assign R24C27_GB10 = R24C27_GBO0;
assign R24C28_GB10 = R24C27_GBO0;
assign R25C26_GB10 = R25C27_GBO0;
assign R25C27_GB10 = R25C27_GBO0;
assign R25C28_GB10 = R25C27_GBO0;
assign R26C26_GB10 = R26C27_GBO0;
assign R26C27_GB10 = R26C27_GBO0;
assign R26C28_GB10 = R26C27_GBO0;
assign R27C26_GB10 = R27C27_GBO0;
assign R27C27_GB10 = R27C27_GBO0;
assign R27C28_GB10 = R27C27_GBO0;
assign R11C2_GB20 = R11C2_GBO0;
assign R11C3_GB20 = R11C2_GBO0;
assign R11C4_GB20 = R11C2_GBO0;
assign R12C2_GB20 = R12C2_GBO0;
assign R12C3_GB20 = R12C2_GBO0;
assign R12C4_GB20 = R12C2_GBO0;
assign R13C2_GB20 = R13C2_GBO0;
assign R13C3_GB20 = R13C2_GBO0;
assign R13C4_GB20 = R13C2_GBO0;
assign R14C2_GB20 = R14C2_GBO0;
assign R14C3_GB20 = R14C2_GBO0;
assign R14C4_GB20 = R14C2_GBO0;
assign R15C2_GB20 = R15C2_GBO0;
assign R15C3_GB20 = R15C2_GBO0;
assign R15C4_GB20 = R15C2_GBO0;
assign R16C2_GB20 = R16C2_GBO0;
assign R16C3_GB20 = R16C2_GBO0;
assign R16C4_GB20 = R16C2_GBO0;
assign R17C2_GB20 = R17C2_GBO0;
assign R17C3_GB20 = R17C2_GBO0;
assign R17C4_GB20 = R17C2_GBO0;
assign R18C2_GB20 = R18C2_GBO0;
assign R18C3_GB20 = R18C2_GBO0;
assign R18C4_GB20 = R18C2_GBO0;
assign R20C2_GB20 = R20C2_GBO0;
assign R20C3_GB20 = R20C2_GBO0;
assign R20C4_GB20 = R20C2_GBO0;
assign R21C2_GB20 = R21C2_GBO0;
assign R21C3_GB20 = R21C2_GBO0;
assign R21C4_GB20 = R21C2_GBO0;
assign R22C2_GB20 = R22C2_GBO0;
assign R22C3_GB20 = R22C2_GBO0;
assign R22C4_GB20 = R22C2_GBO0;
assign R23C2_GB20 = R23C2_GBO0;
assign R23C3_GB20 = R23C2_GBO0;
assign R23C4_GB20 = R23C2_GBO0;
assign R24C2_GB20 = R24C2_GBO0;
assign R24C3_GB20 = R24C2_GBO0;
assign R24C4_GB20 = R24C2_GBO0;
assign R25C2_GB20 = R25C2_GBO0;
assign R25C3_GB20 = R25C2_GBO0;
assign R25C4_GB20 = R25C2_GBO0;
assign R26C2_GB20 = R26C2_GBO0;
assign R26C3_GB20 = R26C2_GBO0;
assign R26C4_GB20 = R26C2_GBO0;
assign R27C2_GB20 = R27C2_GBO0;
assign R27C3_GB20 = R27C2_GBO0;
assign R27C4_GB20 = R27C2_GBO0;
assign R11C5_GB20 = R11C6_GBO0;
assign R11C6_GB20 = R11C6_GBO0;
assign R11C7_GB20 = R11C6_GBO0;
assign R11C8_GB20 = R11C6_GBO0;
assign R12C5_GB20 = R12C6_GBO0;
assign R12C6_GB20 = R12C6_GBO0;
assign R12C7_GB20 = R12C6_GBO0;
assign R12C8_GB20 = R12C6_GBO0;
assign R13C5_GB20 = R13C6_GBO0;
assign R13C6_GB20 = R13C6_GBO0;
assign R13C7_GB20 = R13C6_GBO0;
assign R13C8_GB20 = R13C6_GBO0;
assign R14C5_GB20 = R14C6_GBO0;
assign R14C6_GB20 = R14C6_GBO0;
assign R14C7_GB20 = R14C6_GBO0;
assign R14C8_GB20 = R14C6_GBO0;
assign R15C5_GB20 = R15C6_GBO0;
assign R15C6_GB20 = R15C6_GBO0;
assign R15C7_GB20 = R15C6_GBO0;
assign R15C8_GB20 = R15C6_GBO0;
assign R16C5_GB20 = R16C6_GBO0;
assign R16C6_GB20 = R16C6_GBO0;
assign R16C7_GB20 = R16C6_GBO0;
assign R16C8_GB20 = R16C6_GBO0;
assign R17C5_GB20 = R17C6_GBO0;
assign R17C6_GB20 = R17C6_GBO0;
assign R17C7_GB20 = R17C6_GBO0;
assign R17C8_GB20 = R17C6_GBO0;
assign R18C5_GB20 = R18C6_GBO0;
assign R18C6_GB20 = R18C6_GBO0;
assign R18C7_GB20 = R18C6_GBO0;
assign R18C8_GB20 = R18C6_GBO0;
assign R20C5_GB20 = R20C6_GBO0;
assign R20C6_GB20 = R20C6_GBO0;
assign R20C7_GB20 = R20C6_GBO0;
assign R20C8_GB20 = R20C6_GBO0;
assign R21C5_GB20 = R21C6_GBO0;
assign R21C6_GB20 = R21C6_GBO0;
assign R21C7_GB20 = R21C6_GBO0;
assign R21C8_GB20 = R21C6_GBO0;
assign R22C5_GB20 = R22C6_GBO0;
assign R22C6_GB20 = R22C6_GBO0;
assign R22C7_GB20 = R22C6_GBO0;
assign R22C8_GB20 = R22C6_GBO0;
assign R23C5_GB20 = R23C6_GBO0;
assign R23C6_GB20 = R23C6_GBO0;
assign R23C7_GB20 = R23C6_GBO0;
assign R23C8_GB20 = R23C6_GBO0;
assign R24C5_GB20 = R24C6_GBO0;
assign R24C6_GB20 = R24C6_GBO0;
assign R24C7_GB20 = R24C6_GBO0;
assign R24C8_GB20 = R24C6_GBO0;
assign R25C5_GB20 = R25C6_GBO0;
assign R25C6_GB20 = R25C6_GBO0;
assign R25C7_GB20 = R25C6_GBO0;
assign R25C8_GB20 = R25C6_GBO0;
assign R26C5_GB20 = R26C6_GBO0;
assign R26C6_GB20 = R26C6_GBO0;
assign R26C7_GB20 = R26C6_GBO0;
assign R26C8_GB20 = R26C6_GBO0;
assign R27C5_GB20 = R27C6_GBO0;
assign R27C6_GB20 = R27C6_GBO0;
assign R27C7_GB20 = R27C6_GBO0;
assign R27C8_GB20 = R27C6_GBO0;
assign R11C9_GB20 = R11C10_GBO0;
assign R11C10_GB20 = R11C10_GBO0;
assign R11C11_GB20 = R11C10_GBO0;
assign R11C12_GB20 = R11C10_GBO0;
assign R12C9_GB20 = R12C10_GBO0;
assign R12C10_GB20 = R12C10_GBO0;
assign R12C11_GB20 = R12C10_GBO0;
assign R12C12_GB20 = R12C10_GBO0;
assign R13C9_GB20 = R13C10_GBO0;
assign R13C10_GB20 = R13C10_GBO0;
assign R13C11_GB20 = R13C10_GBO0;
assign R13C12_GB20 = R13C10_GBO0;
assign R14C9_GB20 = R14C10_GBO0;
assign R14C10_GB20 = R14C10_GBO0;
assign R14C11_GB20 = R14C10_GBO0;
assign R14C12_GB20 = R14C10_GBO0;
assign R15C9_GB20 = R15C10_GBO0;
assign R15C10_GB20 = R15C10_GBO0;
assign R15C11_GB20 = R15C10_GBO0;
assign R15C12_GB20 = R15C10_GBO0;
assign R16C9_GB20 = R16C10_GBO0;
assign R16C10_GB20 = R16C10_GBO0;
assign R16C11_GB20 = R16C10_GBO0;
assign R16C12_GB20 = R16C10_GBO0;
assign R17C9_GB20 = R17C10_GBO0;
assign R17C10_GB20 = R17C10_GBO0;
assign R17C11_GB20 = R17C10_GBO0;
assign R17C12_GB20 = R17C10_GBO0;
assign R18C9_GB20 = R18C10_GBO0;
assign R18C10_GB20 = R18C10_GBO0;
assign R18C11_GB20 = R18C10_GBO0;
assign R18C12_GB20 = R18C10_GBO0;
assign R20C9_GB20 = R20C10_GBO0;
assign R20C10_GB20 = R20C10_GBO0;
assign R20C11_GB20 = R20C10_GBO0;
assign R20C12_GB20 = R20C10_GBO0;
assign R21C9_GB20 = R21C10_GBO0;
assign R21C10_GB20 = R21C10_GBO0;
assign R21C11_GB20 = R21C10_GBO0;
assign R21C12_GB20 = R21C10_GBO0;
assign R22C9_GB20 = R22C10_GBO0;
assign R22C10_GB20 = R22C10_GBO0;
assign R22C11_GB20 = R22C10_GBO0;
assign R22C12_GB20 = R22C10_GBO0;
assign R23C9_GB20 = R23C10_GBO0;
assign R23C10_GB20 = R23C10_GBO0;
assign R23C11_GB20 = R23C10_GBO0;
assign R23C12_GB20 = R23C10_GBO0;
assign R24C9_GB20 = R24C10_GBO0;
assign R24C10_GB20 = R24C10_GBO0;
assign R24C11_GB20 = R24C10_GBO0;
assign R24C12_GB20 = R24C10_GBO0;
assign R25C9_GB20 = R25C10_GBO0;
assign R25C10_GB20 = R25C10_GBO0;
assign R25C11_GB20 = R25C10_GBO0;
assign R25C12_GB20 = R25C10_GBO0;
assign R26C9_GB20 = R26C10_GBO0;
assign R26C10_GB20 = R26C10_GBO0;
assign R26C11_GB20 = R26C10_GBO0;
assign R26C12_GB20 = R26C10_GBO0;
assign R27C9_GB20 = R27C10_GBO0;
assign R27C10_GB20 = R27C10_GBO0;
assign R27C11_GB20 = R27C10_GBO0;
assign R27C12_GB20 = R27C10_GBO0;
assign R11C13_GB20 = R11C14_GBO0;
assign R11C14_GB20 = R11C14_GBO0;
assign R11C15_GB20 = R11C14_GBO0;
assign R11C16_GB20 = R11C14_GBO0;
assign R12C13_GB20 = R12C14_GBO0;
assign R12C14_GB20 = R12C14_GBO0;
assign R12C15_GB20 = R12C14_GBO0;
assign R12C16_GB20 = R12C14_GBO0;
assign R13C13_GB20 = R13C14_GBO0;
assign R13C14_GB20 = R13C14_GBO0;
assign R13C15_GB20 = R13C14_GBO0;
assign R13C16_GB20 = R13C14_GBO0;
assign R14C13_GB20 = R14C14_GBO0;
assign R14C14_GB20 = R14C14_GBO0;
assign R14C15_GB20 = R14C14_GBO0;
assign R14C16_GB20 = R14C14_GBO0;
assign R15C13_GB20 = R15C14_GBO0;
assign R15C14_GB20 = R15C14_GBO0;
assign R15C15_GB20 = R15C14_GBO0;
assign R15C16_GB20 = R15C14_GBO0;
assign R16C13_GB20 = R16C14_GBO0;
assign R16C14_GB20 = R16C14_GBO0;
assign R16C15_GB20 = R16C14_GBO0;
assign R16C16_GB20 = R16C14_GBO0;
assign R17C13_GB20 = R17C14_GBO0;
assign R17C14_GB20 = R17C14_GBO0;
assign R17C15_GB20 = R17C14_GBO0;
assign R17C16_GB20 = R17C14_GBO0;
assign R18C13_GB20 = R18C14_GBO0;
assign R18C14_GB20 = R18C14_GBO0;
assign R18C15_GB20 = R18C14_GBO0;
assign R18C16_GB20 = R18C14_GBO0;
assign R20C13_GB20 = R20C14_GBO0;
assign R20C14_GB20 = R20C14_GBO0;
assign R20C15_GB20 = R20C14_GBO0;
assign R20C16_GB20 = R20C14_GBO0;
assign R21C13_GB20 = R21C14_GBO0;
assign R21C14_GB20 = R21C14_GBO0;
assign R21C15_GB20 = R21C14_GBO0;
assign R21C16_GB20 = R21C14_GBO0;
assign R22C13_GB20 = R22C14_GBO0;
assign R22C14_GB20 = R22C14_GBO0;
assign R22C15_GB20 = R22C14_GBO0;
assign R22C16_GB20 = R22C14_GBO0;
assign R23C13_GB20 = R23C14_GBO0;
assign R23C14_GB20 = R23C14_GBO0;
assign R23C15_GB20 = R23C14_GBO0;
assign R23C16_GB20 = R23C14_GBO0;
assign R24C13_GB20 = R24C14_GBO0;
assign R24C14_GB20 = R24C14_GBO0;
assign R24C15_GB20 = R24C14_GBO0;
assign R24C16_GB20 = R24C14_GBO0;
assign R25C13_GB20 = R25C14_GBO0;
assign R25C14_GB20 = R25C14_GBO0;
assign R25C15_GB20 = R25C14_GBO0;
assign R25C16_GB20 = R25C14_GBO0;
assign R26C13_GB20 = R26C14_GBO0;
assign R26C14_GB20 = R26C14_GBO0;
assign R26C15_GB20 = R26C14_GBO0;
assign R26C16_GB20 = R26C14_GBO0;
assign R27C13_GB20 = R27C14_GBO0;
assign R27C14_GB20 = R27C14_GBO0;
assign R27C15_GB20 = R27C14_GBO0;
assign R27C16_GB20 = R27C14_GBO0;
assign R11C17_GB20 = R11C18_GBO0;
assign R11C18_GB20 = R11C18_GBO0;
assign R11C19_GB20 = R11C18_GBO0;
assign R11C20_GB20 = R11C18_GBO0;
assign R12C17_GB20 = R12C18_GBO0;
assign R12C18_GB20 = R12C18_GBO0;
assign R12C19_GB20 = R12C18_GBO0;
assign R12C20_GB20 = R12C18_GBO0;
assign R13C17_GB20 = R13C18_GBO0;
assign R13C18_GB20 = R13C18_GBO0;
assign R13C19_GB20 = R13C18_GBO0;
assign R13C20_GB20 = R13C18_GBO0;
assign R14C17_GB20 = R14C18_GBO0;
assign R14C18_GB20 = R14C18_GBO0;
assign R14C19_GB20 = R14C18_GBO0;
assign R14C20_GB20 = R14C18_GBO0;
assign R15C17_GB20 = R15C18_GBO0;
assign R15C18_GB20 = R15C18_GBO0;
assign R15C19_GB20 = R15C18_GBO0;
assign R15C20_GB20 = R15C18_GBO0;
assign R16C17_GB20 = R16C18_GBO0;
assign R16C18_GB20 = R16C18_GBO0;
assign R16C19_GB20 = R16C18_GBO0;
assign R16C20_GB20 = R16C18_GBO0;
assign R17C17_GB20 = R17C18_GBO0;
assign R17C18_GB20 = R17C18_GBO0;
assign R17C19_GB20 = R17C18_GBO0;
assign R17C20_GB20 = R17C18_GBO0;
assign R18C17_GB20 = R18C18_GBO0;
assign R18C18_GB20 = R18C18_GBO0;
assign R18C19_GB20 = R18C18_GBO0;
assign R18C20_GB20 = R18C18_GBO0;
assign R20C17_GB20 = R20C18_GBO0;
assign R20C18_GB20 = R20C18_GBO0;
assign R20C19_GB20 = R20C18_GBO0;
assign R20C20_GB20 = R20C18_GBO0;
assign R21C17_GB20 = R21C18_GBO0;
assign R21C18_GB20 = R21C18_GBO0;
assign R21C19_GB20 = R21C18_GBO0;
assign R21C20_GB20 = R21C18_GBO0;
assign R22C17_GB20 = R22C18_GBO0;
assign R22C18_GB20 = R22C18_GBO0;
assign R22C19_GB20 = R22C18_GBO0;
assign R22C20_GB20 = R22C18_GBO0;
assign R23C17_GB20 = R23C18_GBO0;
assign R23C18_GB20 = R23C18_GBO0;
assign R23C19_GB20 = R23C18_GBO0;
assign R23C20_GB20 = R23C18_GBO0;
assign R24C17_GB20 = R24C18_GBO0;
assign R24C18_GB20 = R24C18_GBO0;
assign R24C19_GB20 = R24C18_GBO0;
assign R24C20_GB20 = R24C18_GBO0;
assign R25C17_GB20 = R25C18_GBO0;
assign R25C18_GB20 = R25C18_GBO0;
assign R25C19_GB20 = R25C18_GBO0;
assign R25C20_GB20 = R25C18_GBO0;
assign R26C17_GB20 = R26C18_GBO0;
assign R26C18_GB20 = R26C18_GBO0;
assign R26C19_GB20 = R26C18_GBO0;
assign R26C20_GB20 = R26C18_GBO0;
assign R27C17_GB20 = R27C18_GBO0;
assign R27C18_GB20 = R27C18_GBO0;
assign R27C19_GB20 = R27C18_GBO0;
assign R27C20_GB20 = R27C18_GBO0;
assign R11C21_GB20 = R11C22_GBO0;
assign R11C22_GB20 = R11C22_GBO0;
assign R11C23_GB20 = R11C22_GBO0;
assign R11C24_GB20 = R11C22_GBO0;
assign R12C21_GB20 = R12C22_GBO0;
assign R12C22_GB20 = R12C22_GBO0;
assign R12C23_GB20 = R12C22_GBO0;
assign R12C24_GB20 = R12C22_GBO0;
assign R13C21_GB20 = R13C22_GBO0;
assign R13C22_GB20 = R13C22_GBO0;
assign R13C23_GB20 = R13C22_GBO0;
assign R13C24_GB20 = R13C22_GBO0;
assign R14C21_GB20 = R14C22_GBO0;
assign R14C22_GB20 = R14C22_GBO0;
assign R14C23_GB20 = R14C22_GBO0;
assign R14C24_GB20 = R14C22_GBO0;
assign R15C21_GB20 = R15C22_GBO0;
assign R15C22_GB20 = R15C22_GBO0;
assign R15C23_GB20 = R15C22_GBO0;
assign R15C24_GB20 = R15C22_GBO0;
assign R16C21_GB20 = R16C22_GBO0;
assign R16C22_GB20 = R16C22_GBO0;
assign R16C23_GB20 = R16C22_GBO0;
assign R16C24_GB20 = R16C22_GBO0;
assign R17C21_GB20 = R17C22_GBO0;
assign R17C22_GB20 = R17C22_GBO0;
assign R17C23_GB20 = R17C22_GBO0;
assign R17C24_GB20 = R17C22_GBO0;
assign R18C21_GB20 = R18C22_GBO0;
assign R18C22_GB20 = R18C22_GBO0;
assign R18C23_GB20 = R18C22_GBO0;
assign R18C24_GB20 = R18C22_GBO0;
assign R20C21_GB20 = R20C22_GBO0;
assign R20C22_GB20 = R20C22_GBO0;
assign R20C23_GB20 = R20C22_GBO0;
assign R20C24_GB20 = R20C22_GBO0;
assign R21C21_GB20 = R21C22_GBO0;
assign R21C22_GB20 = R21C22_GBO0;
assign R21C23_GB20 = R21C22_GBO0;
assign R21C24_GB20 = R21C22_GBO0;
assign R22C21_GB20 = R22C22_GBO0;
assign R22C22_GB20 = R22C22_GBO0;
assign R22C23_GB20 = R22C22_GBO0;
assign R22C24_GB20 = R22C22_GBO0;
assign R23C21_GB20 = R23C22_GBO0;
assign R23C22_GB20 = R23C22_GBO0;
assign R23C23_GB20 = R23C22_GBO0;
assign R23C24_GB20 = R23C22_GBO0;
assign R24C21_GB20 = R24C22_GBO0;
assign R24C22_GB20 = R24C22_GBO0;
assign R24C23_GB20 = R24C22_GBO0;
assign R24C24_GB20 = R24C22_GBO0;
assign R25C21_GB20 = R25C22_GBO0;
assign R25C22_GB20 = R25C22_GBO0;
assign R25C23_GB20 = R25C22_GBO0;
assign R25C24_GB20 = R25C22_GBO0;
assign R26C21_GB20 = R26C22_GBO0;
assign R26C22_GB20 = R26C22_GBO0;
assign R26C23_GB20 = R26C22_GBO0;
assign R26C24_GB20 = R26C22_GBO0;
assign R27C21_GB20 = R27C22_GBO0;
assign R27C22_GB20 = R27C22_GBO0;
assign R27C23_GB20 = R27C22_GBO0;
assign R27C24_GB20 = R27C22_GBO0;
assign R11C25_GB20 = R11C26_GBO0;
assign R11C26_GB20 = R11C26_GBO0;
assign R11C27_GB20 = R11C26_GBO0;
assign R11C28_GB20 = R11C26_GBO0;
assign R12C25_GB20 = R12C26_GBO0;
assign R12C26_GB20 = R12C26_GBO0;
assign R12C27_GB20 = R12C26_GBO0;
assign R12C28_GB20 = R12C26_GBO0;
assign R13C25_GB20 = R13C26_GBO0;
assign R13C26_GB20 = R13C26_GBO0;
assign R13C27_GB20 = R13C26_GBO0;
assign R13C28_GB20 = R13C26_GBO0;
assign R14C25_GB20 = R14C26_GBO0;
assign R14C26_GB20 = R14C26_GBO0;
assign R14C27_GB20 = R14C26_GBO0;
assign R14C28_GB20 = R14C26_GBO0;
assign R15C25_GB20 = R15C26_GBO0;
assign R15C26_GB20 = R15C26_GBO0;
assign R15C27_GB20 = R15C26_GBO0;
assign R15C28_GB20 = R15C26_GBO0;
assign R16C25_GB20 = R16C26_GBO0;
assign R16C26_GB20 = R16C26_GBO0;
assign R16C27_GB20 = R16C26_GBO0;
assign R16C28_GB20 = R16C26_GBO0;
assign R17C25_GB20 = R17C26_GBO0;
assign R17C26_GB20 = R17C26_GBO0;
assign R17C27_GB20 = R17C26_GBO0;
assign R17C28_GB20 = R17C26_GBO0;
assign R18C25_GB20 = R18C26_GBO0;
assign R18C26_GB20 = R18C26_GBO0;
assign R18C27_GB20 = R18C26_GBO0;
assign R18C28_GB20 = R18C26_GBO0;
assign R20C25_GB20 = R20C26_GBO0;
assign R20C26_GB20 = R20C26_GBO0;
assign R20C27_GB20 = R20C26_GBO0;
assign R20C28_GB20 = R20C26_GBO0;
assign R21C25_GB20 = R21C26_GBO0;
assign R21C26_GB20 = R21C26_GBO0;
assign R21C27_GB20 = R21C26_GBO0;
assign R21C28_GB20 = R21C26_GBO0;
assign R22C25_GB20 = R22C26_GBO0;
assign R22C26_GB20 = R22C26_GBO0;
assign R22C27_GB20 = R22C26_GBO0;
assign R22C28_GB20 = R22C26_GBO0;
assign R23C25_GB20 = R23C26_GBO0;
assign R23C26_GB20 = R23C26_GBO0;
assign R23C27_GB20 = R23C26_GBO0;
assign R23C28_GB20 = R23C26_GBO0;
assign R24C25_GB20 = R24C26_GBO0;
assign R24C26_GB20 = R24C26_GBO0;
assign R24C27_GB20 = R24C26_GBO0;
assign R24C28_GB20 = R24C26_GBO0;
assign R25C25_GB20 = R25C26_GBO0;
assign R25C26_GB20 = R25C26_GBO0;
assign R25C27_GB20 = R25C26_GBO0;
assign R25C28_GB20 = R25C26_GBO0;
assign R26C25_GB20 = R26C26_GBO0;
assign R26C26_GB20 = R26C26_GBO0;
assign R26C27_GB20 = R26C26_GBO0;
assign R26C28_GB20 = R26C26_GBO0;
assign R27C25_GB20 = R27C26_GBO0;
assign R27C26_GB20 = R27C26_GBO0;
assign R27C27_GB20 = R27C26_GBO0;
assign R27C28_GB20 = R27C26_GBO0;
assign R11C2_GB30 = R11C1_GBO0;
assign R11C3_GB30 = R11C1_GBO0;
assign R12C2_GB30 = R12C1_GBO0;
assign R12C3_GB30 = R12C1_GBO0;
assign R13C2_GB30 = R13C1_GBO0;
assign R13C3_GB30 = R13C1_GBO0;
assign R14C2_GB30 = R14C1_GBO0;
assign R14C3_GB30 = R14C1_GBO0;
assign R15C2_GB30 = R15C1_GBO0;
assign R15C3_GB30 = R15C1_GBO0;
assign R16C2_GB30 = R16C1_GBO0;
assign R16C3_GB30 = R16C1_GBO0;
assign R17C2_GB30 = R17C1_GBO0;
assign R17C3_GB30 = R17C1_GBO0;
assign R18C2_GB30 = R18C1_GBO0;
assign R18C3_GB30 = R18C1_GBO0;
assign R20C2_GB30 = R20C1_GBO0;
assign R20C3_GB30 = R20C1_GBO0;
assign R21C2_GB30 = R21C1_GBO0;
assign R21C3_GB30 = R21C1_GBO0;
assign R22C2_GB30 = R22C1_GBO0;
assign R22C3_GB30 = R22C1_GBO0;
assign R23C2_GB30 = R23C1_GBO0;
assign R23C3_GB30 = R23C1_GBO0;
assign R24C2_GB30 = R24C1_GBO0;
assign R24C3_GB30 = R24C1_GBO0;
assign R25C2_GB30 = R25C1_GBO0;
assign R25C3_GB30 = R25C1_GBO0;
assign R26C2_GB30 = R26C1_GBO0;
assign R26C3_GB30 = R26C1_GBO0;
assign R27C2_GB30 = R27C1_GBO0;
assign R27C3_GB30 = R27C1_GBO0;
assign R11C4_GB30 = R11C5_GBO0;
assign R11C5_GB30 = R11C5_GBO0;
assign R11C6_GB30 = R11C5_GBO0;
assign R11C7_GB30 = R11C5_GBO0;
assign R12C4_GB30 = R12C5_GBO0;
assign R12C5_GB30 = R12C5_GBO0;
assign R12C6_GB30 = R12C5_GBO0;
assign R12C7_GB30 = R12C5_GBO0;
assign R13C4_GB30 = R13C5_GBO0;
assign R13C5_GB30 = R13C5_GBO0;
assign R13C6_GB30 = R13C5_GBO0;
assign R13C7_GB30 = R13C5_GBO0;
assign R14C4_GB30 = R14C5_GBO0;
assign R14C5_GB30 = R14C5_GBO0;
assign R14C6_GB30 = R14C5_GBO0;
assign R14C7_GB30 = R14C5_GBO0;
assign R15C4_GB30 = R15C5_GBO0;
assign R15C5_GB30 = R15C5_GBO0;
assign R15C6_GB30 = R15C5_GBO0;
assign R15C7_GB30 = R15C5_GBO0;
assign R16C4_GB30 = R16C5_GBO0;
assign R16C5_GB30 = R16C5_GBO0;
assign R16C6_GB30 = R16C5_GBO0;
assign R16C7_GB30 = R16C5_GBO0;
assign R17C4_GB30 = R17C5_GBO0;
assign R17C5_GB30 = R17C5_GBO0;
assign R17C6_GB30 = R17C5_GBO0;
assign R17C7_GB30 = R17C5_GBO0;
assign R18C4_GB30 = R18C5_GBO0;
assign R18C5_GB30 = R18C5_GBO0;
assign R18C6_GB30 = R18C5_GBO0;
assign R18C7_GB30 = R18C5_GBO0;
assign R20C4_GB30 = R20C5_GBO0;
assign R20C5_GB30 = R20C5_GBO0;
assign R20C6_GB30 = R20C5_GBO0;
assign R20C7_GB30 = R20C5_GBO0;
assign R21C4_GB30 = R21C5_GBO0;
assign R21C5_GB30 = R21C5_GBO0;
assign R21C6_GB30 = R21C5_GBO0;
assign R21C7_GB30 = R21C5_GBO0;
assign R22C4_GB30 = R22C5_GBO0;
assign R22C5_GB30 = R22C5_GBO0;
assign R22C6_GB30 = R22C5_GBO0;
assign R22C7_GB30 = R22C5_GBO0;
assign R23C4_GB30 = R23C5_GBO0;
assign R23C5_GB30 = R23C5_GBO0;
assign R23C6_GB30 = R23C5_GBO0;
assign R23C7_GB30 = R23C5_GBO0;
assign R24C4_GB30 = R24C5_GBO0;
assign R24C5_GB30 = R24C5_GBO0;
assign R24C6_GB30 = R24C5_GBO0;
assign R24C7_GB30 = R24C5_GBO0;
assign R25C4_GB30 = R25C5_GBO0;
assign R25C5_GB30 = R25C5_GBO0;
assign R25C6_GB30 = R25C5_GBO0;
assign R25C7_GB30 = R25C5_GBO0;
assign R26C4_GB30 = R26C5_GBO0;
assign R26C5_GB30 = R26C5_GBO0;
assign R26C6_GB30 = R26C5_GBO0;
assign R26C7_GB30 = R26C5_GBO0;
assign R27C4_GB30 = R27C5_GBO0;
assign R27C5_GB30 = R27C5_GBO0;
assign R27C6_GB30 = R27C5_GBO0;
assign R27C7_GB30 = R27C5_GBO0;
assign R11C9_GB30 = R11C9_GBO0;
assign R11C10_GB30 = R11C9_GBO0;
assign R11C11_GB30 = R11C9_GBO0;
assign R11C8_GB30 = R11C9_GBO0;
assign R12C9_GB30 = R12C9_GBO0;
assign R12C10_GB30 = R12C9_GBO0;
assign R12C11_GB30 = R12C9_GBO0;
assign R12C8_GB30 = R12C9_GBO0;
assign R13C9_GB30 = R13C9_GBO0;
assign R13C10_GB30 = R13C9_GBO0;
assign R13C11_GB30 = R13C9_GBO0;
assign R13C8_GB30 = R13C9_GBO0;
assign R14C9_GB30 = R14C9_GBO0;
assign R14C10_GB30 = R14C9_GBO0;
assign R14C11_GB30 = R14C9_GBO0;
assign R14C8_GB30 = R14C9_GBO0;
assign R15C9_GB30 = R15C9_GBO0;
assign R15C10_GB30 = R15C9_GBO0;
assign R15C11_GB30 = R15C9_GBO0;
assign R15C8_GB30 = R15C9_GBO0;
assign R16C9_GB30 = R16C9_GBO0;
assign R16C10_GB30 = R16C9_GBO0;
assign R16C11_GB30 = R16C9_GBO0;
assign R16C8_GB30 = R16C9_GBO0;
assign R17C9_GB30 = R17C9_GBO0;
assign R17C10_GB30 = R17C9_GBO0;
assign R17C11_GB30 = R17C9_GBO0;
assign R17C8_GB30 = R17C9_GBO0;
assign R18C9_GB30 = R18C9_GBO0;
assign R18C10_GB30 = R18C9_GBO0;
assign R18C11_GB30 = R18C9_GBO0;
assign R18C8_GB30 = R18C9_GBO0;
assign R20C9_GB30 = R20C9_GBO0;
assign R20C10_GB30 = R20C9_GBO0;
assign R20C11_GB30 = R20C9_GBO0;
assign R20C8_GB30 = R20C9_GBO0;
assign R21C9_GB30 = R21C9_GBO0;
assign R21C10_GB30 = R21C9_GBO0;
assign R21C11_GB30 = R21C9_GBO0;
assign R21C8_GB30 = R21C9_GBO0;
assign R22C9_GB30 = R22C9_GBO0;
assign R22C10_GB30 = R22C9_GBO0;
assign R22C11_GB30 = R22C9_GBO0;
assign R22C8_GB30 = R22C9_GBO0;
assign R23C9_GB30 = R23C9_GBO0;
assign R23C10_GB30 = R23C9_GBO0;
assign R23C11_GB30 = R23C9_GBO0;
assign R23C8_GB30 = R23C9_GBO0;
assign R24C9_GB30 = R24C9_GBO0;
assign R24C10_GB30 = R24C9_GBO0;
assign R24C11_GB30 = R24C9_GBO0;
assign R24C8_GB30 = R24C9_GBO0;
assign R25C9_GB30 = R25C9_GBO0;
assign R25C10_GB30 = R25C9_GBO0;
assign R25C11_GB30 = R25C9_GBO0;
assign R25C8_GB30 = R25C9_GBO0;
assign R26C9_GB30 = R26C9_GBO0;
assign R26C10_GB30 = R26C9_GBO0;
assign R26C11_GB30 = R26C9_GBO0;
assign R26C8_GB30 = R26C9_GBO0;
assign R27C9_GB30 = R27C9_GBO0;
assign R27C10_GB30 = R27C9_GBO0;
assign R27C11_GB30 = R27C9_GBO0;
assign R27C8_GB30 = R27C9_GBO0;
assign R11C12_GB30 = R11C13_GBO0;
assign R11C13_GB30 = R11C13_GBO0;
assign R11C14_GB30 = R11C13_GBO0;
assign R11C15_GB30 = R11C13_GBO0;
assign R12C12_GB30 = R12C13_GBO0;
assign R12C13_GB30 = R12C13_GBO0;
assign R12C14_GB30 = R12C13_GBO0;
assign R12C15_GB30 = R12C13_GBO0;
assign R13C12_GB30 = R13C13_GBO0;
assign R13C13_GB30 = R13C13_GBO0;
assign R13C14_GB30 = R13C13_GBO0;
assign R13C15_GB30 = R13C13_GBO0;
assign R14C12_GB30 = R14C13_GBO0;
assign R14C13_GB30 = R14C13_GBO0;
assign R14C14_GB30 = R14C13_GBO0;
assign R14C15_GB30 = R14C13_GBO0;
assign R15C12_GB30 = R15C13_GBO0;
assign R15C13_GB30 = R15C13_GBO0;
assign R15C14_GB30 = R15C13_GBO0;
assign R15C15_GB30 = R15C13_GBO0;
assign R16C12_GB30 = R16C13_GBO0;
assign R16C13_GB30 = R16C13_GBO0;
assign R16C14_GB30 = R16C13_GBO0;
assign R16C15_GB30 = R16C13_GBO0;
assign R17C12_GB30 = R17C13_GBO0;
assign R17C13_GB30 = R17C13_GBO0;
assign R17C14_GB30 = R17C13_GBO0;
assign R17C15_GB30 = R17C13_GBO0;
assign R18C12_GB30 = R18C13_GBO0;
assign R18C13_GB30 = R18C13_GBO0;
assign R18C14_GB30 = R18C13_GBO0;
assign R18C15_GB30 = R18C13_GBO0;
assign R20C12_GB30 = R20C13_GBO0;
assign R20C13_GB30 = R20C13_GBO0;
assign R20C14_GB30 = R20C13_GBO0;
assign R20C15_GB30 = R20C13_GBO0;
assign R21C12_GB30 = R21C13_GBO0;
assign R21C13_GB30 = R21C13_GBO0;
assign R21C14_GB30 = R21C13_GBO0;
assign R21C15_GB30 = R21C13_GBO0;
assign R22C12_GB30 = R22C13_GBO0;
assign R22C13_GB30 = R22C13_GBO0;
assign R22C14_GB30 = R22C13_GBO0;
assign R22C15_GB30 = R22C13_GBO0;
assign R23C12_GB30 = R23C13_GBO0;
assign R23C13_GB30 = R23C13_GBO0;
assign R23C14_GB30 = R23C13_GBO0;
assign R23C15_GB30 = R23C13_GBO0;
assign R24C12_GB30 = R24C13_GBO0;
assign R24C13_GB30 = R24C13_GBO0;
assign R24C14_GB30 = R24C13_GBO0;
assign R24C15_GB30 = R24C13_GBO0;
assign R25C12_GB30 = R25C13_GBO0;
assign R25C13_GB30 = R25C13_GBO0;
assign R25C14_GB30 = R25C13_GBO0;
assign R25C15_GB30 = R25C13_GBO0;
assign R26C12_GB30 = R26C13_GBO0;
assign R26C13_GB30 = R26C13_GBO0;
assign R26C14_GB30 = R26C13_GBO0;
assign R26C15_GB30 = R26C13_GBO0;
assign R27C12_GB30 = R27C13_GBO0;
assign R27C13_GB30 = R27C13_GBO0;
assign R27C14_GB30 = R27C13_GBO0;
assign R27C15_GB30 = R27C13_GBO0;
assign R11C17_GB30 = R11C17_GBO0;
assign R11C18_GB30 = R11C17_GBO0;
assign R11C19_GB30 = R11C17_GBO0;
assign R11C16_GB30 = R11C17_GBO0;
assign R12C17_GB30 = R12C17_GBO0;
assign R12C18_GB30 = R12C17_GBO0;
assign R12C19_GB30 = R12C17_GBO0;
assign R12C16_GB30 = R12C17_GBO0;
assign R13C17_GB30 = R13C17_GBO0;
assign R13C18_GB30 = R13C17_GBO0;
assign R13C19_GB30 = R13C17_GBO0;
assign R13C16_GB30 = R13C17_GBO0;
assign R14C17_GB30 = R14C17_GBO0;
assign R14C18_GB30 = R14C17_GBO0;
assign R14C19_GB30 = R14C17_GBO0;
assign R14C16_GB30 = R14C17_GBO0;
assign R15C17_GB30 = R15C17_GBO0;
assign R15C18_GB30 = R15C17_GBO0;
assign R15C19_GB30 = R15C17_GBO0;
assign R15C16_GB30 = R15C17_GBO0;
assign R16C17_GB30 = R16C17_GBO0;
assign R16C18_GB30 = R16C17_GBO0;
assign R16C19_GB30 = R16C17_GBO0;
assign R16C16_GB30 = R16C17_GBO0;
assign R17C17_GB30 = R17C17_GBO0;
assign R17C18_GB30 = R17C17_GBO0;
assign R17C19_GB30 = R17C17_GBO0;
assign R17C16_GB30 = R17C17_GBO0;
assign R18C17_GB30 = R18C17_GBO0;
assign R18C18_GB30 = R18C17_GBO0;
assign R18C19_GB30 = R18C17_GBO0;
assign R18C16_GB30 = R18C17_GBO0;
assign R20C17_GB30 = R20C17_GBO0;
assign R20C18_GB30 = R20C17_GBO0;
assign R20C19_GB30 = R20C17_GBO0;
assign R20C16_GB30 = R20C17_GBO0;
assign R21C17_GB30 = R21C17_GBO0;
assign R21C18_GB30 = R21C17_GBO0;
assign R21C19_GB30 = R21C17_GBO0;
assign R21C16_GB30 = R21C17_GBO0;
assign R22C17_GB30 = R22C17_GBO0;
assign R22C18_GB30 = R22C17_GBO0;
assign R22C19_GB30 = R22C17_GBO0;
assign R22C16_GB30 = R22C17_GBO0;
assign R23C17_GB30 = R23C17_GBO0;
assign R23C18_GB30 = R23C17_GBO0;
assign R23C19_GB30 = R23C17_GBO0;
assign R23C16_GB30 = R23C17_GBO0;
assign R24C17_GB30 = R24C17_GBO0;
assign R24C18_GB30 = R24C17_GBO0;
assign R24C19_GB30 = R24C17_GBO0;
assign R24C16_GB30 = R24C17_GBO0;
assign R25C17_GB30 = R25C17_GBO0;
assign R25C18_GB30 = R25C17_GBO0;
assign R25C19_GB30 = R25C17_GBO0;
assign R25C16_GB30 = R25C17_GBO0;
assign R26C17_GB30 = R26C17_GBO0;
assign R26C18_GB30 = R26C17_GBO0;
assign R26C19_GB30 = R26C17_GBO0;
assign R26C16_GB30 = R26C17_GBO0;
assign R27C17_GB30 = R27C17_GBO0;
assign R27C18_GB30 = R27C17_GBO0;
assign R27C19_GB30 = R27C17_GBO0;
assign R27C16_GB30 = R27C17_GBO0;
assign R11C20_GB30 = R11C21_GBO0;
assign R11C21_GB30 = R11C21_GBO0;
assign R11C22_GB30 = R11C21_GBO0;
assign R11C23_GB30 = R11C21_GBO0;
assign R12C20_GB30 = R12C21_GBO0;
assign R12C21_GB30 = R12C21_GBO0;
assign R12C22_GB30 = R12C21_GBO0;
assign R12C23_GB30 = R12C21_GBO0;
assign R13C20_GB30 = R13C21_GBO0;
assign R13C21_GB30 = R13C21_GBO0;
assign R13C22_GB30 = R13C21_GBO0;
assign R13C23_GB30 = R13C21_GBO0;
assign R14C20_GB30 = R14C21_GBO0;
assign R14C21_GB30 = R14C21_GBO0;
assign R14C22_GB30 = R14C21_GBO0;
assign R14C23_GB30 = R14C21_GBO0;
assign R15C20_GB30 = R15C21_GBO0;
assign R15C21_GB30 = R15C21_GBO0;
assign R15C22_GB30 = R15C21_GBO0;
assign R15C23_GB30 = R15C21_GBO0;
assign R16C20_GB30 = R16C21_GBO0;
assign R16C21_GB30 = R16C21_GBO0;
assign R16C22_GB30 = R16C21_GBO0;
assign R16C23_GB30 = R16C21_GBO0;
assign R17C20_GB30 = R17C21_GBO0;
assign R17C21_GB30 = R17C21_GBO0;
assign R17C22_GB30 = R17C21_GBO0;
assign R17C23_GB30 = R17C21_GBO0;
assign R18C20_GB30 = R18C21_GBO0;
assign R18C21_GB30 = R18C21_GBO0;
assign R18C22_GB30 = R18C21_GBO0;
assign R18C23_GB30 = R18C21_GBO0;
assign R20C20_GB30 = R20C21_GBO0;
assign R20C21_GB30 = R20C21_GBO0;
assign R20C22_GB30 = R20C21_GBO0;
assign R20C23_GB30 = R20C21_GBO0;
assign R21C20_GB30 = R21C21_GBO0;
assign R21C21_GB30 = R21C21_GBO0;
assign R21C22_GB30 = R21C21_GBO0;
assign R21C23_GB30 = R21C21_GBO0;
assign R22C20_GB30 = R22C21_GBO0;
assign R22C21_GB30 = R22C21_GBO0;
assign R22C22_GB30 = R22C21_GBO0;
assign R22C23_GB30 = R22C21_GBO0;
assign R23C20_GB30 = R23C21_GBO0;
assign R23C21_GB30 = R23C21_GBO0;
assign R23C22_GB30 = R23C21_GBO0;
assign R23C23_GB30 = R23C21_GBO0;
assign R24C20_GB30 = R24C21_GBO0;
assign R24C21_GB30 = R24C21_GBO0;
assign R24C22_GB30 = R24C21_GBO0;
assign R24C23_GB30 = R24C21_GBO0;
assign R25C20_GB30 = R25C21_GBO0;
assign R25C21_GB30 = R25C21_GBO0;
assign R25C22_GB30 = R25C21_GBO0;
assign R25C23_GB30 = R25C21_GBO0;
assign R26C20_GB30 = R26C21_GBO0;
assign R26C21_GB30 = R26C21_GBO0;
assign R26C22_GB30 = R26C21_GBO0;
assign R26C23_GB30 = R26C21_GBO0;
assign R27C20_GB30 = R27C21_GBO0;
assign R27C21_GB30 = R27C21_GBO0;
assign R27C22_GB30 = R27C21_GBO0;
assign R27C23_GB30 = R27C21_GBO0;
assign R11C24_GB30 = R11C25_GBO0;
assign R11C25_GB30 = R11C25_GBO0;
assign R11C26_GB30 = R11C25_GBO0;
assign R11C27_GB30 = R11C25_GBO0;
assign R11C28_GB30 = R11C25_GBO0;
assign R12C24_GB30 = R12C25_GBO0;
assign R12C25_GB30 = R12C25_GBO0;
assign R12C26_GB30 = R12C25_GBO0;
assign R12C27_GB30 = R12C25_GBO0;
assign R12C28_GB30 = R12C25_GBO0;
assign R13C24_GB30 = R13C25_GBO0;
assign R13C25_GB30 = R13C25_GBO0;
assign R13C26_GB30 = R13C25_GBO0;
assign R13C27_GB30 = R13C25_GBO0;
assign R13C28_GB30 = R13C25_GBO0;
assign R14C24_GB30 = R14C25_GBO0;
assign R14C25_GB30 = R14C25_GBO0;
assign R14C26_GB30 = R14C25_GBO0;
assign R14C27_GB30 = R14C25_GBO0;
assign R14C28_GB30 = R14C25_GBO0;
assign R15C24_GB30 = R15C25_GBO0;
assign R15C25_GB30 = R15C25_GBO0;
assign R15C26_GB30 = R15C25_GBO0;
assign R15C27_GB30 = R15C25_GBO0;
assign R15C28_GB30 = R15C25_GBO0;
assign R16C24_GB30 = R16C25_GBO0;
assign R16C25_GB30 = R16C25_GBO0;
assign R16C26_GB30 = R16C25_GBO0;
assign R16C27_GB30 = R16C25_GBO0;
assign R16C28_GB30 = R16C25_GBO0;
assign R17C24_GB30 = R17C25_GBO0;
assign R17C25_GB30 = R17C25_GBO0;
assign R17C26_GB30 = R17C25_GBO0;
assign R17C27_GB30 = R17C25_GBO0;
assign R17C28_GB30 = R17C25_GBO0;
assign R18C24_GB30 = R18C25_GBO0;
assign R18C25_GB30 = R18C25_GBO0;
assign R18C26_GB30 = R18C25_GBO0;
assign R18C27_GB30 = R18C25_GBO0;
assign R18C28_GB30 = R18C25_GBO0;
assign R20C24_GB30 = R20C25_GBO0;
assign R20C25_GB30 = R20C25_GBO0;
assign R20C26_GB30 = R20C25_GBO0;
assign R20C27_GB30 = R20C25_GBO0;
assign R20C28_GB30 = R20C25_GBO0;
assign R21C24_GB30 = R21C25_GBO0;
assign R21C25_GB30 = R21C25_GBO0;
assign R21C26_GB30 = R21C25_GBO0;
assign R21C27_GB30 = R21C25_GBO0;
assign R21C28_GB30 = R21C25_GBO0;
assign R22C24_GB30 = R22C25_GBO0;
assign R22C25_GB30 = R22C25_GBO0;
assign R22C26_GB30 = R22C25_GBO0;
assign R22C27_GB30 = R22C25_GBO0;
assign R22C28_GB30 = R22C25_GBO0;
assign R23C24_GB30 = R23C25_GBO0;
assign R23C25_GB30 = R23C25_GBO0;
assign R23C26_GB30 = R23C25_GBO0;
assign R23C27_GB30 = R23C25_GBO0;
assign R23C28_GB30 = R23C25_GBO0;
assign R24C24_GB30 = R24C25_GBO0;
assign R24C25_GB30 = R24C25_GBO0;
assign R24C26_GB30 = R24C25_GBO0;
assign R24C27_GB30 = R24C25_GBO0;
assign R24C28_GB30 = R24C25_GBO0;
assign R25C24_GB30 = R25C25_GBO0;
assign R25C25_GB30 = R25C25_GBO0;
assign R25C26_GB30 = R25C25_GBO0;
assign R25C27_GB30 = R25C25_GBO0;
assign R25C28_GB30 = R25C25_GBO0;
assign R26C24_GB30 = R26C25_GBO0;
assign R26C25_GB30 = R26C25_GBO0;
assign R26C26_GB30 = R26C25_GBO0;
assign R26C27_GB30 = R26C25_GBO0;
assign R26C28_GB30 = R26C25_GBO0;
assign R27C24_GB30 = R27C25_GBO0;
assign R27C25_GB30 = R27C25_GBO0;
assign R27C26_GB30 = R27C25_GBO0;
assign R27C27_GB30 = R27C25_GBO0;
assign R27C28_GB30 = R27C25_GBO0;
assign R11C2_GB40 = R11C4_GBO1;
assign R11C3_GB40 = R11C4_GBO1;
assign R11C4_GB40 = R11C4_GBO1;
assign R11C5_GB40 = R11C4_GBO1;
assign R11C6_GB40 = R11C4_GBO1;
assign R12C2_GB40 = R12C4_GBO1;
assign R12C3_GB40 = R12C4_GBO1;
assign R12C4_GB40 = R12C4_GBO1;
assign R12C5_GB40 = R12C4_GBO1;
assign R12C6_GB40 = R12C4_GBO1;
assign R13C2_GB40 = R13C4_GBO1;
assign R13C3_GB40 = R13C4_GBO1;
assign R13C4_GB40 = R13C4_GBO1;
assign R13C5_GB40 = R13C4_GBO1;
assign R13C6_GB40 = R13C4_GBO1;
assign R14C2_GB40 = R14C4_GBO1;
assign R14C3_GB40 = R14C4_GBO1;
assign R14C4_GB40 = R14C4_GBO1;
assign R14C5_GB40 = R14C4_GBO1;
assign R14C6_GB40 = R14C4_GBO1;
assign R15C2_GB40 = R15C4_GBO1;
assign R15C3_GB40 = R15C4_GBO1;
assign R15C4_GB40 = R15C4_GBO1;
assign R15C5_GB40 = R15C4_GBO1;
assign R15C6_GB40 = R15C4_GBO1;
assign R16C2_GB40 = R16C4_GBO1;
assign R16C3_GB40 = R16C4_GBO1;
assign R16C4_GB40 = R16C4_GBO1;
assign R16C5_GB40 = R16C4_GBO1;
assign R16C6_GB40 = R16C4_GBO1;
assign R17C2_GB40 = R17C4_GBO1;
assign R17C3_GB40 = R17C4_GBO1;
assign R17C4_GB40 = R17C4_GBO1;
assign R17C5_GB40 = R17C4_GBO1;
assign R17C6_GB40 = R17C4_GBO1;
assign R18C2_GB40 = R18C4_GBO1;
assign R18C3_GB40 = R18C4_GBO1;
assign R18C4_GB40 = R18C4_GBO1;
assign R18C5_GB40 = R18C4_GBO1;
assign R18C6_GB40 = R18C4_GBO1;
assign R20C2_GB40 = R20C4_GBO1;
assign R20C3_GB40 = R20C4_GBO1;
assign R20C4_GB40 = R20C4_GBO1;
assign R20C5_GB40 = R20C4_GBO1;
assign R20C6_GB40 = R20C4_GBO1;
assign R21C2_GB40 = R21C4_GBO1;
assign R21C3_GB40 = R21C4_GBO1;
assign R21C4_GB40 = R21C4_GBO1;
assign R21C5_GB40 = R21C4_GBO1;
assign R21C6_GB40 = R21C4_GBO1;
assign R22C2_GB40 = R22C4_GBO1;
assign R22C3_GB40 = R22C4_GBO1;
assign R22C4_GB40 = R22C4_GBO1;
assign R22C5_GB40 = R22C4_GBO1;
assign R22C6_GB40 = R22C4_GBO1;
assign R23C2_GB40 = R23C4_GBO1;
assign R23C3_GB40 = R23C4_GBO1;
assign R23C4_GB40 = R23C4_GBO1;
assign R23C5_GB40 = R23C4_GBO1;
assign R23C6_GB40 = R23C4_GBO1;
assign R24C2_GB40 = R24C4_GBO1;
assign R24C3_GB40 = R24C4_GBO1;
assign R24C4_GB40 = R24C4_GBO1;
assign R24C5_GB40 = R24C4_GBO1;
assign R24C6_GB40 = R24C4_GBO1;
assign R25C2_GB40 = R25C4_GBO1;
assign R25C3_GB40 = R25C4_GBO1;
assign R25C4_GB40 = R25C4_GBO1;
assign R25C5_GB40 = R25C4_GBO1;
assign R25C6_GB40 = R25C4_GBO1;
assign R26C2_GB40 = R26C4_GBO1;
assign R26C3_GB40 = R26C4_GBO1;
assign R26C4_GB40 = R26C4_GBO1;
assign R26C5_GB40 = R26C4_GBO1;
assign R26C6_GB40 = R26C4_GBO1;
assign R27C2_GB40 = R27C4_GBO1;
assign R27C3_GB40 = R27C4_GBO1;
assign R27C4_GB40 = R27C4_GBO1;
assign R27C5_GB40 = R27C4_GBO1;
assign R27C6_GB40 = R27C4_GBO1;
assign R11C9_GB40 = R11C8_GBO1;
assign R11C10_GB40 = R11C8_GBO1;
assign R11C7_GB40 = R11C8_GBO1;
assign R11C8_GB40 = R11C8_GBO1;
assign R12C9_GB40 = R12C8_GBO1;
assign R12C10_GB40 = R12C8_GBO1;
assign R12C7_GB40 = R12C8_GBO1;
assign R12C8_GB40 = R12C8_GBO1;
assign R13C9_GB40 = R13C8_GBO1;
assign R13C10_GB40 = R13C8_GBO1;
assign R13C7_GB40 = R13C8_GBO1;
assign R13C8_GB40 = R13C8_GBO1;
assign R14C9_GB40 = R14C8_GBO1;
assign R14C10_GB40 = R14C8_GBO1;
assign R14C7_GB40 = R14C8_GBO1;
assign R14C8_GB40 = R14C8_GBO1;
assign R15C9_GB40 = R15C8_GBO1;
assign R15C10_GB40 = R15C8_GBO1;
assign R15C7_GB40 = R15C8_GBO1;
assign R15C8_GB40 = R15C8_GBO1;
assign R16C9_GB40 = R16C8_GBO1;
assign R16C10_GB40 = R16C8_GBO1;
assign R16C7_GB40 = R16C8_GBO1;
assign R16C8_GB40 = R16C8_GBO1;
assign R17C9_GB40 = R17C8_GBO1;
assign R17C10_GB40 = R17C8_GBO1;
assign R17C7_GB40 = R17C8_GBO1;
assign R17C8_GB40 = R17C8_GBO1;
assign R18C9_GB40 = R18C8_GBO1;
assign R18C10_GB40 = R18C8_GBO1;
assign R18C7_GB40 = R18C8_GBO1;
assign R18C8_GB40 = R18C8_GBO1;
assign R20C9_GB40 = R20C8_GBO1;
assign R20C10_GB40 = R20C8_GBO1;
assign R20C7_GB40 = R20C8_GBO1;
assign R20C8_GB40 = R20C8_GBO1;
assign R21C9_GB40 = R21C8_GBO1;
assign R21C10_GB40 = R21C8_GBO1;
assign R21C7_GB40 = R21C8_GBO1;
assign R21C8_GB40 = R21C8_GBO1;
assign R22C9_GB40 = R22C8_GBO1;
assign R22C10_GB40 = R22C8_GBO1;
assign R22C7_GB40 = R22C8_GBO1;
assign R22C8_GB40 = R22C8_GBO1;
assign R23C9_GB40 = R23C8_GBO1;
assign R23C10_GB40 = R23C8_GBO1;
assign R23C7_GB40 = R23C8_GBO1;
assign R23C8_GB40 = R23C8_GBO1;
assign R24C9_GB40 = R24C8_GBO1;
assign R24C10_GB40 = R24C8_GBO1;
assign R24C7_GB40 = R24C8_GBO1;
assign R24C8_GB40 = R24C8_GBO1;
assign R25C9_GB40 = R25C8_GBO1;
assign R25C10_GB40 = R25C8_GBO1;
assign R25C7_GB40 = R25C8_GBO1;
assign R25C8_GB40 = R25C8_GBO1;
assign R26C9_GB40 = R26C8_GBO1;
assign R26C10_GB40 = R26C8_GBO1;
assign R26C7_GB40 = R26C8_GBO1;
assign R26C8_GB40 = R26C8_GBO1;
assign R27C9_GB40 = R27C8_GBO1;
assign R27C10_GB40 = R27C8_GBO1;
assign R27C7_GB40 = R27C8_GBO1;
assign R27C8_GB40 = R27C8_GBO1;
assign R11C11_GB40 = R11C12_GBO1;
assign R11C12_GB40 = R11C12_GBO1;
assign R11C13_GB40 = R11C12_GBO1;
assign R11C14_GB40 = R11C12_GBO1;
assign R12C11_GB40 = R12C12_GBO1;
assign R12C12_GB40 = R12C12_GBO1;
assign R12C13_GB40 = R12C12_GBO1;
assign R12C14_GB40 = R12C12_GBO1;
assign R13C11_GB40 = R13C12_GBO1;
assign R13C12_GB40 = R13C12_GBO1;
assign R13C13_GB40 = R13C12_GBO1;
assign R13C14_GB40 = R13C12_GBO1;
assign R14C11_GB40 = R14C12_GBO1;
assign R14C12_GB40 = R14C12_GBO1;
assign R14C13_GB40 = R14C12_GBO1;
assign R14C14_GB40 = R14C12_GBO1;
assign R15C11_GB40 = R15C12_GBO1;
assign R15C12_GB40 = R15C12_GBO1;
assign R15C13_GB40 = R15C12_GBO1;
assign R15C14_GB40 = R15C12_GBO1;
assign R16C11_GB40 = R16C12_GBO1;
assign R16C12_GB40 = R16C12_GBO1;
assign R16C13_GB40 = R16C12_GBO1;
assign R16C14_GB40 = R16C12_GBO1;
assign R17C11_GB40 = R17C12_GBO1;
assign R17C12_GB40 = R17C12_GBO1;
assign R17C13_GB40 = R17C12_GBO1;
assign R17C14_GB40 = R17C12_GBO1;
assign R18C11_GB40 = R18C12_GBO1;
assign R18C12_GB40 = R18C12_GBO1;
assign R18C13_GB40 = R18C12_GBO1;
assign R18C14_GB40 = R18C12_GBO1;
assign R20C11_GB40 = R20C12_GBO1;
assign R20C12_GB40 = R20C12_GBO1;
assign R20C13_GB40 = R20C12_GBO1;
assign R20C14_GB40 = R20C12_GBO1;
assign R21C11_GB40 = R21C12_GBO1;
assign R21C12_GB40 = R21C12_GBO1;
assign R21C13_GB40 = R21C12_GBO1;
assign R21C14_GB40 = R21C12_GBO1;
assign R22C11_GB40 = R22C12_GBO1;
assign R22C12_GB40 = R22C12_GBO1;
assign R22C13_GB40 = R22C12_GBO1;
assign R22C14_GB40 = R22C12_GBO1;
assign R23C11_GB40 = R23C12_GBO1;
assign R23C12_GB40 = R23C12_GBO1;
assign R23C13_GB40 = R23C12_GBO1;
assign R23C14_GB40 = R23C12_GBO1;
assign R24C11_GB40 = R24C12_GBO1;
assign R24C12_GB40 = R24C12_GBO1;
assign R24C13_GB40 = R24C12_GBO1;
assign R24C14_GB40 = R24C12_GBO1;
assign R25C11_GB40 = R25C12_GBO1;
assign R25C12_GB40 = R25C12_GBO1;
assign R25C13_GB40 = R25C12_GBO1;
assign R25C14_GB40 = R25C12_GBO1;
assign R26C11_GB40 = R26C12_GBO1;
assign R26C12_GB40 = R26C12_GBO1;
assign R26C13_GB40 = R26C12_GBO1;
assign R26C14_GB40 = R26C12_GBO1;
assign R27C11_GB40 = R27C12_GBO1;
assign R27C12_GB40 = R27C12_GBO1;
assign R27C13_GB40 = R27C12_GBO1;
assign R27C14_GB40 = R27C12_GBO1;
assign R11C17_GB40 = R11C16_GBO1;
assign R11C18_GB40 = R11C16_GBO1;
assign R11C15_GB40 = R11C16_GBO1;
assign R11C16_GB40 = R11C16_GBO1;
assign R12C17_GB40 = R12C16_GBO1;
assign R12C18_GB40 = R12C16_GBO1;
assign R12C15_GB40 = R12C16_GBO1;
assign R12C16_GB40 = R12C16_GBO1;
assign R13C17_GB40 = R13C16_GBO1;
assign R13C18_GB40 = R13C16_GBO1;
assign R13C15_GB40 = R13C16_GBO1;
assign R13C16_GB40 = R13C16_GBO1;
assign R14C17_GB40 = R14C16_GBO1;
assign R14C18_GB40 = R14C16_GBO1;
assign R14C15_GB40 = R14C16_GBO1;
assign R14C16_GB40 = R14C16_GBO1;
assign R15C17_GB40 = R15C16_GBO1;
assign R15C18_GB40 = R15C16_GBO1;
assign R15C15_GB40 = R15C16_GBO1;
assign R15C16_GB40 = R15C16_GBO1;
assign R16C17_GB40 = R16C16_GBO1;
assign R16C18_GB40 = R16C16_GBO1;
assign R16C15_GB40 = R16C16_GBO1;
assign R16C16_GB40 = R16C16_GBO1;
assign R17C17_GB40 = R17C16_GBO1;
assign R17C18_GB40 = R17C16_GBO1;
assign R17C15_GB40 = R17C16_GBO1;
assign R17C16_GB40 = R17C16_GBO1;
assign R18C17_GB40 = R18C16_GBO1;
assign R18C18_GB40 = R18C16_GBO1;
assign R18C15_GB40 = R18C16_GBO1;
assign R18C16_GB40 = R18C16_GBO1;
assign R20C17_GB40 = R20C16_GBO1;
assign R20C18_GB40 = R20C16_GBO1;
assign R20C15_GB40 = R20C16_GBO1;
assign R20C16_GB40 = R20C16_GBO1;
assign R21C17_GB40 = R21C16_GBO1;
assign R21C18_GB40 = R21C16_GBO1;
assign R21C15_GB40 = R21C16_GBO1;
assign R21C16_GB40 = R21C16_GBO1;
assign R22C17_GB40 = R22C16_GBO1;
assign R22C18_GB40 = R22C16_GBO1;
assign R22C15_GB40 = R22C16_GBO1;
assign R22C16_GB40 = R22C16_GBO1;
assign R23C17_GB40 = R23C16_GBO1;
assign R23C18_GB40 = R23C16_GBO1;
assign R23C15_GB40 = R23C16_GBO1;
assign R23C16_GB40 = R23C16_GBO1;
assign R24C17_GB40 = R24C16_GBO1;
assign R24C18_GB40 = R24C16_GBO1;
assign R24C15_GB40 = R24C16_GBO1;
assign R24C16_GB40 = R24C16_GBO1;
assign R25C17_GB40 = R25C16_GBO1;
assign R25C18_GB40 = R25C16_GBO1;
assign R25C15_GB40 = R25C16_GBO1;
assign R25C16_GB40 = R25C16_GBO1;
assign R26C17_GB40 = R26C16_GBO1;
assign R26C18_GB40 = R26C16_GBO1;
assign R26C15_GB40 = R26C16_GBO1;
assign R26C16_GB40 = R26C16_GBO1;
assign R27C17_GB40 = R27C16_GBO1;
assign R27C18_GB40 = R27C16_GBO1;
assign R27C15_GB40 = R27C16_GBO1;
assign R27C16_GB40 = R27C16_GBO1;
assign R11C19_GB40 = R11C20_GBO1;
assign R11C20_GB40 = R11C20_GBO1;
assign R11C21_GB40 = R11C20_GBO1;
assign R11C22_GB40 = R11C20_GBO1;
assign R12C19_GB40 = R12C20_GBO1;
assign R12C20_GB40 = R12C20_GBO1;
assign R12C21_GB40 = R12C20_GBO1;
assign R12C22_GB40 = R12C20_GBO1;
assign R13C19_GB40 = R13C20_GBO1;
assign R13C20_GB40 = R13C20_GBO1;
assign R13C21_GB40 = R13C20_GBO1;
assign R13C22_GB40 = R13C20_GBO1;
assign R14C19_GB40 = R14C20_GBO1;
assign R14C20_GB40 = R14C20_GBO1;
assign R14C21_GB40 = R14C20_GBO1;
assign R14C22_GB40 = R14C20_GBO1;
assign R15C19_GB40 = R15C20_GBO1;
assign R15C20_GB40 = R15C20_GBO1;
assign R15C21_GB40 = R15C20_GBO1;
assign R15C22_GB40 = R15C20_GBO1;
assign R16C19_GB40 = R16C20_GBO1;
assign R16C20_GB40 = R16C20_GBO1;
assign R16C21_GB40 = R16C20_GBO1;
assign R16C22_GB40 = R16C20_GBO1;
assign R17C19_GB40 = R17C20_GBO1;
assign R17C20_GB40 = R17C20_GBO1;
assign R17C21_GB40 = R17C20_GBO1;
assign R17C22_GB40 = R17C20_GBO1;
assign R18C19_GB40 = R18C20_GBO1;
assign R18C20_GB40 = R18C20_GBO1;
assign R18C21_GB40 = R18C20_GBO1;
assign R18C22_GB40 = R18C20_GBO1;
assign R20C19_GB40 = R20C20_GBO1;
assign R20C20_GB40 = R20C20_GBO1;
assign R20C21_GB40 = R20C20_GBO1;
assign R20C22_GB40 = R20C20_GBO1;
assign R21C19_GB40 = R21C20_GBO1;
assign R21C20_GB40 = R21C20_GBO1;
assign R21C21_GB40 = R21C20_GBO1;
assign R21C22_GB40 = R21C20_GBO1;
assign R22C19_GB40 = R22C20_GBO1;
assign R22C20_GB40 = R22C20_GBO1;
assign R22C21_GB40 = R22C20_GBO1;
assign R22C22_GB40 = R22C20_GBO1;
assign R23C19_GB40 = R23C20_GBO1;
assign R23C20_GB40 = R23C20_GBO1;
assign R23C21_GB40 = R23C20_GBO1;
assign R23C22_GB40 = R23C20_GBO1;
assign R24C19_GB40 = R24C20_GBO1;
assign R24C20_GB40 = R24C20_GBO1;
assign R24C21_GB40 = R24C20_GBO1;
assign R24C22_GB40 = R24C20_GBO1;
assign R25C19_GB40 = R25C20_GBO1;
assign R25C20_GB40 = R25C20_GBO1;
assign R25C21_GB40 = R25C20_GBO1;
assign R25C22_GB40 = R25C20_GBO1;
assign R26C19_GB40 = R26C20_GBO1;
assign R26C20_GB40 = R26C20_GBO1;
assign R26C21_GB40 = R26C20_GBO1;
assign R26C22_GB40 = R26C20_GBO1;
assign R27C19_GB40 = R27C20_GBO1;
assign R27C20_GB40 = R27C20_GBO1;
assign R27C21_GB40 = R27C20_GBO1;
assign R27C22_GB40 = R27C20_GBO1;
assign R11C23_GB40 = R11C24_GBO1;
assign R11C24_GB40 = R11C24_GBO1;
assign R11C25_GB40 = R11C24_GBO1;
assign R11C26_GB40 = R11C24_GBO1;
assign R11C27_GB40 = R11C24_GBO1;
assign R11C28_GB40 = R11C24_GBO1;
assign R12C23_GB40 = R12C24_GBO1;
assign R12C24_GB40 = R12C24_GBO1;
assign R12C25_GB40 = R12C24_GBO1;
assign R12C26_GB40 = R12C24_GBO1;
assign R12C27_GB40 = R12C24_GBO1;
assign R12C28_GB40 = R12C24_GBO1;
assign R13C23_GB40 = R13C24_GBO1;
assign R13C24_GB40 = R13C24_GBO1;
assign R13C25_GB40 = R13C24_GBO1;
assign R13C26_GB40 = R13C24_GBO1;
assign R13C27_GB40 = R13C24_GBO1;
assign R13C28_GB40 = R13C24_GBO1;
assign R14C23_GB40 = R14C24_GBO1;
assign R14C24_GB40 = R14C24_GBO1;
assign R14C25_GB40 = R14C24_GBO1;
assign R14C26_GB40 = R14C24_GBO1;
assign R14C27_GB40 = R14C24_GBO1;
assign R14C28_GB40 = R14C24_GBO1;
assign R15C23_GB40 = R15C24_GBO1;
assign R15C24_GB40 = R15C24_GBO1;
assign R15C25_GB40 = R15C24_GBO1;
assign R15C26_GB40 = R15C24_GBO1;
assign R15C27_GB40 = R15C24_GBO1;
assign R15C28_GB40 = R15C24_GBO1;
assign R16C23_GB40 = R16C24_GBO1;
assign R16C24_GB40 = R16C24_GBO1;
assign R16C25_GB40 = R16C24_GBO1;
assign R16C26_GB40 = R16C24_GBO1;
assign R16C27_GB40 = R16C24_GBO1;
assign R16C28_GB40 = R16C24_GBO1;
assign R17C23_GB40 = R17C24_GBO1;
assign R17C24_GB40 = R17C24_GBO1;
assign R17C25_GB40 = R17C24_GBO1;
assign R17C26_GB40 = R17C24_GBO1;
assign R17C27_GB40 = R17C24_GBO1;
assign R17C28_GB40 = R17C24_GBO1;
assign R18C23_GB40 = R18C24_GBO1;
assign R18C24_GB40 = R18C24_GBO1;
assign R18C25_GB40 = R18C24_GBO1;
assign R18C26_GB40 = R18C24_GBO1;
assign R18C27_GB40 = R18C24_GBO1;
assign R18C28_GB40 = R18C24_GBO1;
assign R20C23_GB40 = R20C24_GBO1;
assign R20C24_GB40 = R20C24_GBO1;
assign R20C25_GB40 = R20C24_GBO1;
assign R20C26_GB40 = R20C24_GBO1;
assign R20C27_GB40 = R20C24_GBO1;
assign R20C28_GB40 = R20C24_GBO1;
assign R21C23_GB40 = R21C24_GBO1;
assign R21C24_GB40 = R21C24_GBO1;
assign R21C25_GB40 = R21C24_GBO1;
assign R21C26_GB40 = R21C24_GBO1;
assign R21C27_GB40 = R21C24_GBO1;
assign R21C28_GB40 = R21C24_GBO1;
assign R22C23_GB40 = R22C24_GBO1;
assign R22C24_GB40 = R22C24_GBO1;
assign R22C25_GB40 = R22C24_GBO1;
assign R22C26_GB40 = R22C24_GBO1;
assign R22C27_GB40 = R22C24_GBO1;
assign R22C28_GB40 = R22C24_GBO1;
assign R23C23_GB40 = R23C24_GBO1;
assign R23C24_GB40 = R23C24_GBO1;
assign R23C25_GB40 = R23C24_GBO1;
assign R23C26_GB40 = R23C24_GBO1;
assign R23C27_GB40 = R23C24_GBO1;
assign R23C28_GB40 = R23C24_GBO1;
assign R24C23_GB40 = R24C24_GBO1;
assign R24C24_GB40 = R24C24_GBO1;
assign R24C25_GB40 = R24C24_GBO1;
assign R24C26_GB40 = R24C24_GBO1;
assign R24C27_GB40 = R24C24_GBO1;
assign R24C28_GB40 = R24C24_GBO1;
assign R25C23_GB40 = R25C24_GBO1;
assign R25C24_GB40 = R25C24_GBO1;
assign R25C25_GB40 = R25C24_GBO1;
assign R25C26_GB40 = R25C24_GBO1;
assign R25C27_GB40 = R25C24_GBO1;
assign R25C28_GB40 = R25C24_GBO1;
assign R26C23_GB40 = R26C24_GBO1;
assign R26C24_GB40 = R26C24_GBO1;
assign R26C25_GB40 = R26C24_GBO1;
assign R26C26_GB40 = R26C24_GBO1;
assign R26C27_GB40 = R26C24_GBO1;
assign R26C28_GB40 = R26C24_GBO1;
assign R27C23_GB40 = R27C24_GBO1;
assign R27C24_GB40 = R27C24_GBO1;
assign R27C25_GB40 = R27C24_GBO1;
assign R27C26_GB40 = R27C24_GBO1;
assign R27C27_GB40 = R27C24_GBO1;
assign R27C28_GB40 = R27C24_GBO1;
assign R11C2_GB50 = R11C3_GBO1;
assign R11C3_GB50 = R11C3_GBO1;
assign R11C4_GB50 = R11C3_GBO1;
assign R11C5_GB50 = R11C3_GBO1;
assign R12C2_GB50 = R12C3_GBO1;
assign R12C3_GB50 = R12C3_GBO1;
assign R12C4_GB50 = R12C3_GBO1;
assign R12C5_GB50 = R12C3_GBO1;
assign R13C2_GB50 = R13C3_GBO1;
assign R13C3_GB50 = R13C3_GBO1;
assign R13C4_GB50 = R13C3_GBO1;
assign R13C5_GB50 = R13C3_GBO1;
assign R14C2_GB50 = R14C3_GBO1;
assign R14C3_GB50 = R14C3_GBO1;
assign R14C4_GB50 = R14C3_GBO1;
assign R14C5_GB50 = R14C3_GBO1;
assign R15C2_GB50 = R15C3_GBO1;
assign R15C3_GB50 = R15C3_GBO1;
assign R15C4_GB50 = R15C3_GBO1;
assign R15C5_GB50 = R15C3_GBO1;
assign R16C2_GB50 = R16C3_GBO1;
assign R16C3_GB50 = R16C3_GBO1;
assign R16C4_GB50 = R16C3_GBO1;
assign R16C5_GB50 = R16C3_GBO1;
assign R17C2_GB50 = R17C3_GBO1;
assign R17C3_GB50 = R17C3_GBO1;
assign R17C4_GB50 = R17C3_GBO1;
assign R17C5_GB50 = R17C3_GBO1;
assign R18C2_GB50 = R18C3_GBO1;
assign R18C3_GB50 = R18C3_GBO1;
assign R18C4_GB50 = R18C3_GBO1;
assign R18C5_GB50 = R18C3_GBO1;
assign R20C2_GB50 = R20C3_GBO1;
assign R20C3_GB50 = R20C3_GBO1;
assign R20C4_GB50 = R20C3_GBO1;
assign R20C5_GB50 = R20C3_GBO1;
assign R21C2_GB50 = R21C3_GBO1;
assign R21C3_GB50 = R21C3_GBO1;
assign R21C4_GB50 = R21C3_GBO1;
assign R21C5_GB50 = R21C3_GBO1;
assign R22C2_GB50 = R22C3_GBO1;
assign R22C3_GB50 = R22C3_GBO1;
assign R22C4_GB50 = R22C3_GBO1;
assign R22C5_GB50 = R22C3_GBO1;
assign R23C2_GB50 = R23C3_GBO1;
assign R23C3_GB50 = R23C3_GBO1;
assign R23C4_GB50 = R23C3_GBO1;
assign R23C5_GB50 = R23C3_GBO1;
assign R24C2_GB50 = R24C3_GBO1;
assign R24C3_GB50 = R24C3_GBO1;
assign R24C4_GB50 = R24C3_GBO1;
assign R24C5_GB50 = R24C3_GBO1;
assign R25C2_GB50 = R25C3_GBO1;
assign R25C3_GB50 = R25C3_GBO1;
assign R25C4_GB50 = R25C3_GBO1;
assign R25C5_GB50 = R25C3_GBO1;
assign R26C2_GB50 = R26C3_GBO1;
assign R26C3_GB50 = R26C3_GBO1;
assign R26C4_GB50 = R26C3_GBO1;
assign R26C5_GB50 = R26C3_GBO1;
assign R27C2_GB50 = R27C3_GBO1;
assign R27C3_GB50 = R27C3_GBO1;
assign R27C4_GB50 = R27C3_GBO1;
assign R27C5_GB50 = R27C3_GBO1;
assign R11C9_GB50 = R11C7_GBO1;
assign R11C6_GB50 = R11C7_GBO1;
assign R11C7_GB50 = R11C7_GBO1;
assign R11C8_GB50 = R11C7_GBO1;
assign R12C9_GB50 = R12C7_GBO1;
assign R12C6_GB50 = R12C7_GBO1;
assign R12C7_GB50 = R12C7_GBO1;
assign R12C8_GB50 = R12C7_GBO1;
assign R13C9_GB50 = R13C7_GBO1;
assign R13C6_GB50 = R13C7_GBO1;
assign R13C7_GB50 = R13C7_GBO1;
assign R13C8_GB50 = R13C7_GBO1;
assign R14C9_GB50 = R14C7_GBO1;
assign R14C6_GB50 = R14C7_GBO1;
assign R14C7_GB50 = R14C7_GBO1;
assign R14C8_GB50 = R14C7_GBO1;
assign R15C9_GB50 = R15C7_GBO1;
assign R15C6_GB50 = R15C7_GBO1;
assign R15C7_GB50 = R15C7_GBO1;
assign R15C8_GB50 = R15C7_GBO1;
assign R16C9_GB50 = R16C7_GBO1;
assign R16C6_GB50 = R16C7_GBO1;
assign R16C7_GB50 = R16C7_GBO1;
assign R16C8_GB50 = R16C7_GBO1;
assign R17C9_GB50 = R17C7_GBO1;
assign R17C6_GB50 = R17C7_GBO1;
assign R17C7_GB50 = R17C7_GBO1;
assign R17C8_GB50 = R17C7_GBO1;
assign R18C9_GB50 = R18C7_GBO1;
assign R18C6_GB50 = R18C7_GBO1;
assign R18C7_GB50 = R18C7_GBO1;
assign R18C8_GB50 = R18C7_GBO1;
assign R20C9_GB50 = R20C7_GBO1;
assign R20C6_GB50 = R20C7_GBO1;
assign R20C7_GB50 = R20C7_GBO1;
assign R20C8_GB50 = R20C7_GBO1;
assign R21C9_GB50 = R21C7_GBO1;
assign R21C6_GB50 = R21C7_GBO1;
assign R21C7_GB50 = R21C7_GBO1;
assign R21C8_GB50 = R21C7_GBO1;
assign R22C9_GB50 = R22C7_GBO1;
assign R22C6_GB50 = R22C7_GBO1;
assign R22C7_GB50 = R22C7_GBO1;
assign R22C8_GB50 = R22C7_GBO1;
assign R23C9_GB50 = R23C7_GBO1;
assign R23C6_GB50 = R23C7_GBO1;
assign R23C7_GB50 = R23C7_GBO1;
assign R23C8_GB50 = R23C7_GBO1;
assign R24C9_GB50 = R24C7_GBO1;
assign R24C6_GB50 = R24C7_GBO1;
assign R24C7_GB50 = R24C7_GBO1;
assign R24C8_GB50 = R24C7_GBO1;
assign R25C9_GB50 = R25C7_GBO1;
assign R25C6_GB50 = R25C7_GBO1;
assign R25C7_GB50 = R25C7_GBO1;
assign R25C8_GB50 = R25C7_GBO1;
assign R26C9_GB50 = R26C7_GBO1;
assign R26C6_GB50 = R26C7_GBO1;
assign R26C7_GB50 = R26C7_GBO1;
assign R26C8_GB50 = R26C7_GBO1;
assign R27C9_GB50 = R27C7_GBO1;
assign R27C6_GB50 = R27C7_GBO1;
assign R27C7_GB50 = R27C7_GBO1;
assign R27C8_GB50 = R27C7_GBO1;
assign R11C10_GB50 = R11C11_GBO1;
assign R11C11_GB50 = R11C11_GBO1;
assign R11C12_GB50 = R11C11_GBO1;
assign R11C13_GB50 = R11C11_GBO1;
assign R12C10_GB50 = R12C11_GBO1;
assign R12C11_GB50 = R12C11_GBO1;
assign R12C12_GB50 = R12C11_GBO1;
assign R12C13_GB50 = R12C11_GBO1;
assign R13C10_GB50 = R13C11_GBO1;
assign R13C11_GB50 = R13C11_GBO1;
assign R13C12_GB50 = R13C11_GBO1;
assign R13C13_GB50 = R13C11_GBO1;
assign R14C10_GB50 = R14C11_GBO1;
assign R14C11_GB50 = R14C11_GBO1;
assign R14C12_GB50 = R14C11_GBO1;
assign R14C13_GB50 = R14C11_GBO1;
assign R15C10_GB50 = R15C11_GBO1;
assign R15C11_GB50 = R15C11_GBO1;
assign R15C12_GB50 = R15C11_GBO1;
assign R15C13_GB50 = R15C11_GBO1;
assign R16C10_GB50 = R16C11_GBO1;
assign R16C11_GB50 = R16C11_GBO1;
assign R16C12_GB50 = R16C11_GBO1;
assign R16C13_GB50 = R16C11_GBO1;
assign R17C10_GB50 = R17C11_GBO1;
assign R17C11_GB50 = R17C11_GBO1;
assign R17C12_GB50 = R17C11_GBO1;
assign R17C13_GB50 = R17C11_GBO1;
assign R18C10_GB50 = R18C11_GBO1;
assign R18C11_GB50 = R18C11_GBO1;
assign R18C12_GB50 = R18C11_GBO1;
assign R18C13_GB50 = R18C11_GBO1;
assign R20C10_GB50 = R20C11_GBO1;
assign R20C11_GB50 = R20C11_GBO1;
assign R20C12_GB50 = R20C11_GBO1;
assign R20C13_GB50 = R20C11_GBO1;
assign R21C10_GB50 = R21C11_GBO1;
assign R21C11_GB50 = R21C11_GBO1;
assign R21C12_GB50 = R21C11_GBO1;
assign R21C13_GB50 = R21C11_GBO1;
assign R22C10_GB50 = R22C11_GBO1;
assign R22C11_GB50 = R22C11_GBO1;
assign R22C12_GB50 = R22C11_GBO1;
assign R22C13_GB50 = R22C11_GBO1;
assign R23C10_GB50 = R23C11_GBO1;
assign R23C11_GB50 = R23C11_GBO1;
assign R23C12_GB50 = R23C11_GBO1;
assign R23C13_GB50 = R23C11_GBO1;
assign R24C10_GB50 = R24C11_GBO1;
assign R24C11_GB50 = R24C11_GBO1;
assign R24C12_GB50 = R24C11_GBO1;
assign R24C13_GB50 = R24C11_GBO1;
assign R25C10_GB50 = R25C11_GBO1;
assign R25C11_GB50 = R25C11_GBO1;
assign R25C12_GB50 = R25C11_GBO1;
assign R25C13_GB50 = R25C11_GBO1;
assign R26C10_GB50 = R26C11_GBO1;
assign R26C11_GB50 = R26C11_GBO1;
assign R26C12_GB50 = R26C11_GBO1;
assign R26C13_GB50 = R26C11_GBO1;
assign R27C10_GB50 = R27C11_GBO1;
assign R27C11_GB50 = R27C11_GBO1;
assign R27C12_GB50 = R27C11_GBO1;
assign R27C13_GB50 = R27C11_GBO1;
assign R11C17_GB50 = R11C15_GBO1;
assign R11C14_GB50 = R11C15_GBO1;
assign R11C15_GB50 = R11C15_GBO1;
assign R11C16_GB50 = R11C15_GBO1;
assign R12C17_GB50 = R12C15_GBO1;
assign R12C14_GB50 = R12C15_GBO1;
assign R12C15_GB50 = R12C15_GBO1;
assign R12C16_GB50 = R12C15_GBO1;
assign R13C17_GB50 = R13C15_GBO1;
assign R13C14_GB50 = R13C15_GBO1;
assign R13C15_GB50 = R13C15_GBO1;
assign R13C16_GB50 = R13C15_GBO1;
assign R14C17_GB50 = R14C15_GBO1;
assign R14C14_GB50 = R14C15_GBO1;
assign R14C15_GB50 = R14C15_GBO1;
assign R14C16_GB50 = R14C15_GBO1;
assign R15C17_GB50 = R15C15_GBO1;
assign R15C14_GB50 = R15C15_GBO1;
assign R15C15_GB50 = R15C15_GBO1;
assign R15C16_GB50 = R15C15_GBO1;
assign R16C17_GB50 = R16C15_GBO1;
assign R16C14_GB50 = R16C15_GBO1;
assign R16C15_GB50 = R16C15_GBO1;
assign R16C16_GB50 = R16C15_GBO1;
assign R17C17_GB50 = R17C15_GBO1;
assign R17C14_GB50 = R17C15_GBO1;
assign R17C15_GB50 = R17C15_GBO1;
assign R17C16_GB50 = R17C15_GBO1;
assign R18C17_GB50 = R18C15_GBO1;
assign R18C14_GB50 = R18C15_GBO1;
assign R18C15_GB50 = R18C15_GBO1;
assign R18C16_GB50 = R18C15_GBO1;
assign R20C17_GB50 = R20C15_GBO1;
assign R20C14_GB50 = R20C15_GBO1;
assign R20C15_GB50 = R20C15_GBO1;
assign R20C16_GB50 = R20C15_GBO1;
assign R21C17_GB50 = R21C15_GBO1;
assign R21C14_GB50 = R21C15_GBO1;
assign R21C15_GB50 = R21C15_GBO1;
assign R21C16_GB50 = R21C15_GBO1;
assign R22C17_GB50 = R22C15_GBO1;
assign R22C14_GB50 = R22C15_GBO1;
assign R22C15_GB50 = R22C15_GBO1;
assign R22C16_GB50 = R22C15_GBO1;
assign R23C17_GB50 = R23C15_GBO1;
assign R23C14_GB50 = R23C15_GBO1;
assign R23C15_GB50 = R23C15_GBO1;
assign R23C16_GB50 = R23C15_GBO1;
assign R24C17_GB50 = R24C15_GBO1;
assign R24C14_GB50 = R24C15_GBO1;
assign R24C15_GB50 = R24C15_GBO1;
assign R24C16_GB50 = R24C15_GBO1;
assign R25C17_GB50 = R25C15_GBO1;
assign R25C14_GB50 = R25C15_GBO1;
assign R25C15_GB50 = R25C15_GBO1;
assign R25C16_GB50 = R25C15_GBO1;
assign R26C17_GB50 = R26C15_GBO1;
assign R26C14_GB50 = R26C15_GBO1;
assign R26C15_GB50 = R26C15_GBO1;
assign R26C16_GB50 = R26C15_GBO1;
assign R27C17_GB50 = R27C15_GBO1;
assign R27C14_GB50 = R27C15_GBO1;
assign R27C15_GB50 = R27C15_GBO1;
assign R27C16_GB50 = R27C15_GBO1;
assign R11C18_GB50 = R11C19_GBO1;
assign R11C19_GB50 = R11C19_GBO1;
assign R11C20_GB50 = R11C19_GBO1;
assign R11C21_GB50 = R11C19_GBO1;
assign R12C18_GB50 = R12C19_GBO1;
assign R12C19_GB50 = R12C19_GBO1;
assign R12C20_GB50 = R12C19_GBO1;
assign R12C21_GB50 = R12C19_GBO1;
assign R13C18_GB50 = R13C19_GBO1;
assign R13C19_GB50 = R13C19_GBO1;
assign R13C20_GB50 = R13C19_GBO1;
assign R13C21_GB50 = R13C19_GBO1;
assign R14C18_GB50 = R14C19_GBO1;
assign R14C19_GB50 = R14C19_GBO1;
assign R14C20_GB50 = R14C19_GBO1;
assign R14C21_GB50 = R14C19_GBO1;
assign R15C18_GB50 = R15C19_GBO1;
assign R15C19_GB50 = R15C19_GBO1;
assign R15C20_GB50 = R15C19_GBO1;
assign R15C21_GB50 = R15C19_GBO1;
assign R16C18_GB50 = R16C19_GBO1;
assign R16C19_GB50 = R16C19_GBO1;
assign R16C20_GB50 = R16C19_GBO1;
assign R16C21_GB50 = R16C19_GBO1;
assign R17C18_GB50 = R17C19_GBO1;
assign R17C19_GB50 = R17C19_GBO1;
assign R17C20_GB50 = R17C19_GBO1;
assign R17C21_GB50 = R17C19_GBO1;
assign R18C18_GB50 = R18C19_GBO1;
assign R18C19_GB50 = R18C19_GBO1;
assign R18C20_GB50 = R18C19_GBO1;
assign R18C21_GB50 = R18C19_GBO1;
assign R20C18_GB50 = R20C19_GBO1;
assign R20C19_GB50 = R20C19_GBO1;
assign R20C20_GB50 = R20C19_GBO1;
assign R20C21_GB50 = R20C19_GBO1;
assign R21C18_GB50 = R21C19_GBO1;
assign R21C19_GB50 = R21C19_GBO1;
assign R21C20_GB50 = R21C19_GBO1;
assign R21C21_GB50 = R21C19_GBO1;
assign R22C18_GB50 = R22C19_GBO1;
assign R22C19_GB50 = R22C19_GBO1;
assign R22C20_GB50 = R22C19_GBO1;
assign R22C21_GB50 = R22C19_GBO1;
assign R23C18_GB50 = R23C19_GBO1;
assign R23C19_GB50 = R23C19_GBO1;
assign R23C20_GB50 = R23C19_GBO1;
assign R23C21_GB50 = R23C19_GBO1;
assign R24C18_GB50 = R24C19_GBO1;
assign R24C19_GB50 = R24C19_GBO1;
assign R24C20_GB50 = R24C19_GBO1;
assign R24C21_GB50 = R24C19_GBO1;
assign R25C18_GB50 = R25C19_GBO1;
assign R25C19_GB50 = R25C19_GBO1;
assign R25C20_GB50 = R25C19_GBO1;
assign R25C21_GB50 = R25C19_GBO1;
assign R26C18_GB50 = R26C19_GBO1;
assign R26C19_GB50 = R26C19_GBO1;
assign R26C20_GB50 = R26C19_GBO1;
assign R26C21_GB50 = R26C19_GBO1;
assign R27C18_GB50 = R27C19_GBO1;
assign R27C19_GB50 = R27C19_GBO1;
assign R27C20_GB50 = R27C19_GBO1;
assign R27C21_GB50 = R27C19_GBO1;
assign R11C25_GB50 = R11C23_GBO1;
assign R11C22_GB50 = R11C23_GBO1;
assign R11C23_GB50 = R11C23_GBO1;
assign R11C24_GB50 = R11C23_GBO1;
assign R12C25_GB50 = R12C23_GBO1;
assign R12C22_GB50 = R12C23_GBO1;
assign R12C23_GB50 = R12C23_GBO1;
assign R12C24_GB50 = R12C23_GBO1;
assign R13C25_GB50 = R13C23_GBO1;
assign R13C22_GB50 = R13C23_GBO1;
assign R13C23_GB50 = R13C23_GBO1;
assign R13C24_GB50 = R13C23_GBO1;
assign R14C25_GB50 = R14C23_GBO1;
assign R14C22_GB50 = R14C23_GBO1;
assign R14C23_GB50 = R14C23_GBO1;
assign R14C24_GB50 = R14C23_GBO1;
assign R15C25_GB50 = R15C23_GBO1;
assign R15C22_GB50 = R15C23_GBO1;
assign R15C23_GB50 = R15C23_GBO1;
assign R15C24_GB50 = R15C23_GBO1;
assign R16C25_GB50 = R16C23_GBO1;
assign R16C22_GB50 = R16C23_GBO1;
assign R16C23_GB50 = R16C23_GBO1;
assign R16C24_GB50 = R16C23_GBO1;
assign R17C25_GB50 = R17C23_GBO1;
assign R17C22_GB50 = R17C23_GBO1;
assign R17C23_GB50 = R17C23_GBO1;
assign R17C24_GB50 = R17C23_GBO1;
assign R18C25_GB50 = R18C23_GBO1;
assign R18C22_GB50 = R18C23_GBO1;
assign R18C23_GB50 = R18C23_GBO1;
assign R18C24_GB50 = R18C23_GBO1;
assign R20C25_GB50 = R20C23_GBO1;
assign R20C22_GB50 = R20C23_GBO1;
assign R20C23_GB50 = R20C23_GBO1;
assign R20C24_GB50 = R20C23_GBO1;
assign R21C25_GB50 = R21C23_GBO1;
assign R21C22_GB50 = R21C23_GBO1;
assign R21C23_GB50 = R21C23_GBO1;
assign R21C24_GB50 = R21C23_GBO1;
assign R22C25_GB50 = R22C23_GBO1;
assign R22C22_GB50 = R22C23_GBO1;
assign R22C23_GB50 = R22C23_GBO1;
assign R22C24_GB50 = R22C23_GBO1;
assign R23C25_GB50 = R23C23_GBO1;
assign R23C22_GB50 = R23C23_GBO1;
assign R23C23_GB50 = R23C23_GBO1;
assign R23C24_GB50 = R23C23_GBO1;
assign R24C25_GB50 = R24C23_GBO1;
assign R24C22_GB50 = R24C23_GBO1;
assign R24C23_GB50 = R24C23_GBO1;
assign R24C24_GB50 = R24C23_GBO1;
assign R25C25_GB50 = R25C23_GBO1;
assign R25C22_GB50 = R25C23_GBO1;
assign R25C23_GB50 = R25C23_GBO1;
assign R25C24_GB50 = R25C23_GBO1;
assign R26C25_GB50 = R26C23_GBO1;
assign R26C22_GB50 = R26C23_GBO1;
assign R26C23_GB50 = R26C23_GBO1;
assign R26C24_GB50 = R26C23_GBO1;
assign R27C25_GB50 = R27C23_GBO1;
assign R27C22_GB50 = R27C23_GBO1;
assign R27C23_GB50 = R27C23_GBO1;
assign R27C24_GB50 = R27C23_GBO1;
assign R11C26_GB50 = R11C27_GBO1;
assign R11C27_GB50 = R11C27_GBO1;
assign R11C28_GB50 = R11C27_GBO1;
assign R12C26_GB50 = R12C27_GBO1;
assign R12C27_GB50 = R12C27_GBO1;
assign R12C28_GB50 = R12C27_GBO1;
assign R13C26_GB50 = R13C27_GBO1;
assign R13C27_GB50 = R13C27_GBO1;
assign R13C28_GB50 = R13C27_GBO1;
assign R14C26_GB50 = R14C27_GBO1;
assign R14C27_GB50 = R14C27_GBO1;
assign R14C28_GB50 = R14C27_GBO1;
assign R15C26_GB50 = R15C27_GBO1;
assign R15C27_GB50 = R15C27_GBO1;
assign R15C28_GB50 = R15C27_GBO1;
assign R16C26_GB50 = R16C27_GBO1;
assign R16C27_GB50 = R16C27_GBO1;
assign R16C28_GB50 = R16C27_GBO1;
assign R17C26_GB50 = R17C27_GBO1;
assign R17C27_GB50 = R17C27_GBO1;
assign R17C28_GB50 = R17C27_GBO1;
assign R18C26_GB50 = R18C27_GBO1;
assign R18C27_GB50 = R18C27_GBO1;
assign R18C28_GB50 = R18C27_GBO1;
assign R20C26_GB50 = R20C27_GBO1;
assign R20C27_GB50 = R20C27_GBO1;
assign R20C28_GB50 = R20C27_GBO1;
assign R21C26_GB50 = R21C27_GBO1;
assign R21C27_GB50 = R21C27_GBO1;
assign R21C28_GB50 = R21C27_GBO1;
assign R22C26_GB50 = R22C27_GBO1;
assign R22C27_GB50 = R22C27_GBO1;
assign R22C28_GB50 = R22C27_GBO1;
assign R23C26_GB50 = R23C27_GBO1;
assign R23C27_GB50 = R23C27_GBO1;
assign R23C28_GB50 = R23C27_GBO1;
assign R24C26_GB50 = R24C27_GBO1;
assign R24C27_GB50 = R24C27_GBO1;
assign R24C28_GB50 = R24C27_GBO1;
assign R25C26_GB50 = R25C27_GBO1;
assign R25C27_GB50 = R25C27_GBO1;
assign R25C28_GB50 = R25C27_GBO1;
assign R26C26_GB50 = R26C27_GBO1;
assign R26C27_GB50 = R26C27_GBO1;
assign R26C28_GB50 = R26C27_GBO1;
assign R27C26_GB50 = R27C27_GBO1;
assign R27C27_GB50 = R27C27_GBO1;
assign R27C28_GB50 = R27C27_GBO1;
assign R11C2_GB60 = R11C2_GBO1;
assign R11C3_GB60 = R11C2_GBO1;
assign R11C4_GB60 = R11C2_GBO1;
assign R12C2_GB60 = R12C2_GBO1;
assign R12C3_GB60 = R12C2_GBO1;
assign R12C4_GB60 = R12C2_GBO1;
assign R13C2_GB60 = R13C2_GBO1;
assign R13C3_GB60 = R13C2_GBO1;
assign R13C4_GB60 = R13C2_GBO1;
assign R14C2_GB60 = R14C2_GBO1;
assign R14C3_GB60 = R14C2_GBO1;
assign R14C4_GB60 = R14C2_GBO1;
assign R15C2_GB60 = R15C2_GBO1;
assign R15C3_GB60 = R15C2_GBO1;
assign R15C4_GB60 = R15C2_GBO1;
assign R16C2_GB60 = R16C2_GBO1;
assign R16C3_GB60 = R16C2_GBO1;
assign R16C4_GB60 = R16C2_GBO1;
assign R17C2_GB60 = R17C2_GBO1;
assign R17C3_GB60 = R17C2_GBO1;
assign R17C4_GB60 = R17C2_GBO1;
assign R18C2_GB60 = R18C2_GBO1;
assign R18C3_GB60 = R18C2_GBO1;
assign R18C4_GB60 = R18C2_GBO1;
assign R20C2_GB60 = R20C2_GBO1;
assign R20C3_GB60 = R20C2_GBO1;
assign R20C4_GB60 = R20C2_GBO1;
assign R21C2_GB60 = R21C2_GBO1;
assign R21C3_GB60 = R21C2_GBO1;
assign R21C4_GB60 = R21C2_GBO1;
assign R22C2_GB60 = R22C2_GBO1;
assign R22C3_GB60 = R22C2_GBO1;
assign R22C4_GB60 = R22C2_GBO1;
assign R23C2_GB60 = R23C2_GBO1;
assign R23C3_GB60 = R23C2_GBO1;
assign R23C4_GB60 = R23C2_GBO1;
assign R24C2_GB60 = R24C2_GBO1;
assign R24C3_GB60 = R24C2_GBO1;
assign R24C4_GB60 = R24C2_GBO1;
assign R25C2_GB60 = R25C2_GBO1;
assign R25C3_GB60 = R25C2_GBO1;
assign R25C4_GB60 = R25C2_GBO1;
assign R26C2_GB60 = R26C2_GBO1;
assign R26C3_GB60 = R26C2_GBO1;
assign R26C4_GB60 = R26C2_GBO1;
assign R27C2_GB60 = R27C2_GBO1;
assign R27C3_GB60 = R27C2_GBO1;
assign R27C4_GB60 = R27C2_GBO1;
assign R11C5_GB60 = R11C6_GBO1;
assign R11C6_GB60 = R11C6_GBO1;
assign R11C7_GB60 = R11C6_GBO1;
assign R11C8_GB60 = R11C6_GBO1;
assign R12C5_GB60 = R12C6_GBO1;
assign R12C6_GB60 = R12C6_GBO1;
assign R12C7_GB60 = R12C6_GBO1;
assign R12C8_GB60 = R12C6_GBO1;
assign R13C5_GB60 = R13C6_GBO1;
assign R13C6_GB60 = R13C6_GBO1;
assign R13C7_GB60 = R13C6_GBO1;
assign R13C8_GB60 = R13C6_GBO1;
assign R14C5_GB60 = R14C6_GBO1;
assign R14C6_GB60 = R14C6_GBO1;
assign R14C7_GB60 = R14C6_GBO1;
assign R14C8_GB60 = R14C6_GBO1;
assign R15C5_GB60 = R15C6_GBO1;
assign R15C6_GB60 = R15C6_GBO1;
assign R15C7_GB60 = R15C6_GBO1;
assign R15C8_GB60 = R15C6_GBO1;
assign R16C5_GB60 = R16C6_GBO1;
assign R16C6_GB60 = R16C6_GBO1;
assign R16C7_GB60 = R16C6_GBO1;
assign R16C8_GB60 = R16C6_GBO1;
assign R17C5_GB60 = R17C6_GBO1;
assign R17C6_GB60 = R17C6_GBO1;
assign R17C7_GB60 = R17C6_GBO1;
assign R17C8_GB60 = R17C6_GBO1;
assign R18C5_GB60 = R18C6_GBO1;
assign R18C6_GB60 = R18C6_GBO1;
assign R18C7_GB60 = R18C6_GBO1;
assign R18C8_GB60 = R18C6_GBO1;
assign R20C5_GB60 = R20C6_GBO1;
assign R20C6_GB60 = R20C6_GBO1;
assign R20C7_GB60 = R20C6_GBO1;
assign R20C8_GB60 = R20C6_GBO1;
assign R21C5_GB60 = R21C6_GBO1;
assign R21C6_GB60 = R21C6_GBO1;
assign R21C7_GB60 = R21C6_GBO1;
assign R21C8_GB60 = R21C6_GBO1;
assign R22C5_GB60 = R22C6_GBO1;
assign R22C6_GB60 = R22C6_GBO1;
assign R22C7_GB60 = R22C6_GBO1;
assign R22C8_GB60 = R22C6_GBO1;
assign R23C5_GB60 = R23C6_GBO1;
assign R23C6_GB60 = R23C6_GBO1;
assign R23C7_GB60 = R23C6_GBO1;
assign R23C8_GB60 = R23C6_GBO1;
assign R24C5_GB60 = R24C6_GBO1;
assign R24C6_GB60 = R24C6_GBO1;
assign R24C7_GB60 = R24C6_GBO1;
assign R24C8_GB60 = R24C6_GBO1;
assign R25C5_GB60 = R25C6_GBO1;
assign R25C6_GB60 = R25C6_GBO1;
assign R25C7_GB60 = R25C6_GBO1;
assign R25C8_GB60 = R25C6_GBO1;
assign R26C5_GB60 = R26C6_GBO1;
assign R26C6_GB60 = R26C6_GBO1;
assign R26C7_GB60 = R26C6_GBO1;
assign R26C8_GB60 = R26C6_GBO1;
assign R27C5_GB60 = R27C6_GBO1;
assign R27C6_GB60 = R27C6_GBO1;
assign R27C7_GB60 = R27C6_GBO1;
assign R27C8_GB60 = R27C6_GBO1;
assign R11C9_GB60 = R11C10_GBO1;
assign R11C10_GB60 = R11C10_GBO1;
assign R11C11_GB60 = R11C10_GBO1;
assign R11C12_GB60 = R11C10_GBO1;
assign R12C9_GB60 = R12C10_GBO1;
assign R12C10_GB60 = R12C10_GBO1;
assign R12C11_GB60 = R12C10_GBO1;
assign R12C12_GB60 = R12C10_GBO1;
assign R13C9_GB60 = R13C10_GBO1;
assign R13C10_GB60 = R13C10_GBO1;
assign R13C11_GB60 = R13C10_GBO1;
assign R13C12_GB60 = R13C10_GBO1;
assign R14C9_GB60 = R14C10_GBO1;
assign R14C10_GB60 = R14C10_GBO1;
assign R14C11_GB60 = R14C10_GBO1;
assign R14C12_GB60 = R14C10_GBO1;
assign R15C9_GB60 = R15C10_GBO1;
assign R15C10_GB60 = R15C10_GBO1;
assign R15C11_GB60 = R15C10_GBO1;
assign R15C12_GB60 = R15C10_GBO1;
assign R16C9_GB60 = R16C10_GBO1;
assign R16C10_GB60 = R16C10_GBO1;
assign R16C11_GB60 = R16C10_GBO1;
assign R16C12_GB60 = R16C10_GBO1;
assign R17C9_GB60 = R17C10_GBO1;
assign R17C10_GB60 = R17C10_GBO1;
assign R17C11_GB60 = R17C10_GBO1;
assign R17C12_GB60 = R17C10_GBO1;
assign R18C9_GB60 = R18C10_GBO1;
assign R18C10_GB60 = R18C10_GBO1;
assign R18C11_GB60 = R18C10_GBO1;
assign R18C12_GB60 = R18C10_GBO1;
assign R20C9_GB60 = R20C10_GBO1;
assign R20C10_GB60 = R20C10_GBO1;
assign R20C11_GB60 = R20C10_GBO1;
assign R20C12_GB60 = R20C10_GBO1;
assign R21C9_GB60 = R21C10_GBO1;
assign R21C10_GB60 = R21C10_GBO1;
assign R21C11_GB60 = R21C10_GBO1;
assign R21C12_GB60 = R21C10_GBO1;
assign R22C9_GB60 = R22C10_GBO1;
assign R22C10_GB60 = R22C10_GBO1;
assign R22C11_GB60 = R22C10_GBO1;
assign R22C12_GB60 = R22C10_GBO1;
assign R23C9_GB60 = R23C10_GBO1;
assign R23C10_GB60 = R23C10_GBO1;
assign R23C11_GB60 = R23C10_GBO1;
assign R23C12_GB60 = R23C10_GBO1;
assign R24C9_GB60 = R24C10_GBO1;
assign R24C10_GB60 = R24C10_GBO1;
assign R24C11_GB60 = R24C10_GBO1;
assign R24C12_GB60 = R24C10_GBO1;
assign R25C9_GB60 = R25C10_GBO1;
assign R25C10_GB60 = R25C10_GBO1;
assign R25C11_GB60 = R25C10_GBO1;
assign R25C12_GB60 = R25C10_GBO1;
assign R26C9_GB60 = R26C10_GBO1;
assign R26C10_GB60 = R26C10_GBO1;
assign R26C11_GB60 = R26C10_GBO1;
assign R26C12_GB60 = R26C10_GBO1;
assign R27C9_GB60 = R27C10_GBO1;
assign R27C10_GB60 = R27C10_GBO1;
assign R27C11_GB60 = R27C10_GBO1;
assign R27C12_GB60 = R27C10_GBO1;
assign R11C13_GB60 = R11C14_GBO1;
assign R11C14_GB60 = R11C14_GBO1;
assign R11C15_GB60 = R11C14_GBO1;
assign R11C16_GB60 = R11C14_GBO1;
assign R12C13_GB60 = R12C14_GBO1;
assign R12C14_GB60 = R12C14_GBO1;
assign R12C15_GB60 = R12C14_GBO1;
assign R12C16_GB60 = R12C14_GBO1;
assign R13C13_GB60 = R13C14_GBO1;
assign R13C14_GB60 = R13C14_GBO1;
assign R13C15_GB60 = R13C14_GBO1;
assign R13C16_GB60 = R13C14_GBO1;
assign R14C13_GB60 = R14C14_GBO1;
assign R14C14_GB60 = R14C14_GBO1;
assign R14C15_GB60 = R14C14_GBO1;
assign R14C16_GB60 = R14C14_GBO1;
assign R15C13_GB60 = R15C14_GBO1;
assign R15C14_GB60 = R15C14_GBO1;
assign R15C15_GB60 = R15C14_GBO1;
assign R15C16_GB60 = R15C14_GBO1;
assign R16C13_GB60 = R16C14_GBO1;
assign R16C14_GB60 = R16C14_GBO1;
assign R16C15_GB60 = R16C14_GBO1;
assign R16C16_GB60 = R16C14_GBO1;
assign R17C13_GB60 = R17C14_GBO1;
assign R17C14_GB60 = R17C14_GBO1;
assign R17C15_GB60 = R17C14_GBO1;
assign R17C16_GB60 = R17C14_GBO1;
assign R18C13_GB60 = R18C14_GBO1;
assign R18C14_GB60 = R18C14_GBO1;
assign R18C15_GB60 = R18C14_GBO1;
assign R18C16_GB60 = R18C14_GBO1;
assign R20C13_GB60 = R20C14_GBO1;
assign R20C14_GB60 = R20C14_GBO1;
assign R20C15_GB60 = R20C14_GBO1;
assign R20C16_GB60 = R20C14_GBO1;
assign R21C13_GB60 = R21C14_GBO1;
assign R21C14_GB60 = R21C14_GBO1;
assign R21C15_GB60 = R21C14_GBO1;
assign R21C16_GB60 = R21C14_GBO1;
assign R22C13_GB60 = R22C14_GBO1;
assign R22C14_GB60 = R22C14_GBO1;
assign R22C15_GB60 = R22C14_GBO1;
assign R22C16_GB60 = R22C14_GBO1;
assign R23C13_GB60 = R23C14_GBO1;
assign R23C14_GB60 = R23C14_GBO1;
assign R23C15_GB60 = R23C14_GBO1;
assign R23C16_GB60 = R23C14_GBO1;
assign R24C13_GB60 = R24C14_GBO1;
assign R24C14_GB60 = R24C14_GBO1;
assign R24C15_GB60 = R24C14_GBO1;
assign R24C16_GB60 = R24C14_GBO1;
assign R25C13_GB60 = R25C14_GBO1;
assign R25C14_GB60 = R25C14_GBO1;
assign R25C15_GB60 = R25C14_GBO1;
assign R25C16_GB60 = R25C14_GBO1;
assign R26C13_GB60 = R26C14_GBO1;
assign R26C14_GB60 = R26C14_GBO1;
assign R26C15_GB60 = R26C14_GBO1;
assign R26C16_GB60 = R26C14_GBO1;
assign R27C13_GB60 = R27C14_GBO1;
assign R27C14_GB60 = R27C14_GBO1;
assign R27C15_GB60 = R27C14_GBO1;
assign R27C16_GB60 = R27C14_GBO1;
assign R11C17_GB60 = R11C18_GBO1;
assign R11C18_GB60 = R11C18_GBO1;
assign R11C19_GB60 = R11C18_GBO1;
assign R11C20_GB60 = R11C18_GBO1;
assign R12C17_GB60 = R12C18_GBO1;
assign R12C18_GB60 = R12C18_GBO1;
assign R12C19_GB60 = R12C18_GBO1;
assign R12C20_GB60 = R12C18_GBO1;
assign R13C17_GB60 = R13C18_GBO1;
assign R13C18_GB60 = R13C18_GBO1;
assign R13C19_GB60 = R13C18_GBO1;
assign R13C20_GB60 = R13C18_GBO1;
assign R14C17_GB60 = R14C18_GBO1;
assign R14C18_GB60 = R14C18_GBO1;
assign R14C19_GB60 = R14C18_GBO1;
assign R14C20_GB60 = R14C18_GBO1;
assign R15C17_GB60 = R15C18_GBO1;
assign R15C18_GB60 = R15C18_GBO1;
assign R15C19_GB60 = R15C18_GBO1;
assign R15C20_GB60 = R15C18_GBO1;
assign R16C17_GB60 = R16C18_GBO1;
assign R16C18_GB60 = R16C18_GBO1;
assign R16C19_GB60 = R16C18_GBO1;
assign R16C20_GB60 = R16C18_GBO1;
assign R17C17_GB60 = R17C18_GBO1;
assign R17C18_GB60 = R17C18_GBO1;
assign R17C19_GB60 = R17C18_GBO1;
assign R17C20_GB60 = R17C18_GBO1;
assign R18C17_GB60 = R18C18_GBO1;
assign R18C18_GB60 = R18C18_GBO1;
assign R18C19_GB60 = R18C18_GBO1;
assign R18C20_GB60 = R18C18_GBO1;
assign R20C17_GB60 = R20C18_GBO1;
assign R20C18_GB60 = R20C18_GBO1;
assign R20C19_GB60 = R20C18_GBO1;
assign R20C20_GB60 = R20C18_GBO1;
assign R21C17_GB60 = R21C18_GBO1;
assign R21C18_GB60 = R21C18_GBO1;
assign R21C19_GB60 = R21C18_GBO1;
assign R21C20_GB60 = R21C18_GBO1;
assign R22C17_GB60 = R22C18_GBO1;
assign R22C18_GB60 = R22C18_GBO1;
assign R22C19_GB60 = R22C18_GBO1;
assign R22C20_GB60 = R22C18_GBO1;
assign R23C17_GB60 = R23C18_GBO1;
assign R23C18_GB60 = R23C18_GBO1;
assign R23C19_GB60 = R23C18_GBO1;
assign R23C20_GB60 = R23C18_GBO1;
assign R24C17_GB60 = R24C18_GBO1;
assign R24C18_GB60 = R24C18_GBO1;
assign R24C19_GB60 = R24C18_GBO1;
assign R24C20_GB60 = R24C18_GBO1;
assign R25C17_GB60 = R25C18_GBO1;
assign R25C18_GB60 = R25C18_GBO1;
assign R25C19_GB60 = R25C18_GBO1;
assign R25C20_GB60 = R25C18_GBO1;
assign R26C17_GB60 = R26C18_GBO1;
assign R26C18_GB60 = R26C18_GBO1;
assign R26C19_GB60 = R26C18_GBO1;
assign R26C20_GB60 = R26C18_GBO1;
assign R27C17_GB60 = R27C18_GBO1;
assign R27C18_GB60 = R27C18_GBO1;
assign R27C19_GB60 = R27C18_GBO1;
assign R27C20_GB60 = R27C18_GBO1;
assign R11C21_GB60 = R11C22_GBO1;
assign R11C22_GB60 = R11C22_GBO1;
assign R11C23_GB60 = R11C22_GBO1;
assign R11C24_GB60 = R11C22_GBO1;
assign R12C21_GB60 = R12C22_GBO1;
assign R12C22_GB60 = R12C22_GBO1;
assign R12C23_GB60 = R12C22_GBO1;
assign R12C24_GB60 = R12C22_GBO1;
assign R13C21_GB60 = R13C22_GBO1;
assign R13C22_GB60 = R13C22_GBO1;
assign R13C23_GB60 = R13C22_GBO1;
assign R13C24_GB60 = R13C22_GBO1;
assign R14C21_GB60 = R14C22_GBO1;
assign R14C22_GB60 = R14C22_GBO1;
assign R14C23_GB60 = R14C22_GBO1;
assign R14C24_GB60 = R14C22_GBO1;
assign R15C21_GB60 = R15C22_GBO1;
assign R15C22_GB60 = R15C22_GBO1;
assign R15C23_GB60 = R15C22_GBO1;
assign R15C24_GB60 = R15C22_GBO1;
assign R16C21_GB60 = R16C22_GBO1;
assign R16C22_GB60 = R16C22_GBO1;
assign R16C23_GB60 = R16C22_GBO1;
assign R16C24_GB60 = R16C22_GBO1;
assign R17C21_GB60 = R17C22_GBO1;
assign R17C22_GB60 = R17C22_GBO1;
assign R17C23_GB60 = R17C22_GBO1;
assign R17C24_GB60 = R17C22_GBO1;
assign R18C21_GB60 = R18C22_GBO1;
assign R18C22_GB60 = R18C22_GBO1;
assign R18C23_GB60 = R18C22_GBO1;
assign R18C24_GB60 = R18C22_GBO1;
assign R20C21_GB60 = R20C22_GBO1;
assign R20C22_GB60 = R20C22_GBO1;
assign R20C23_GB60 = R20C22_GBO1;
assign R20C24_GB60 = R20C22_GBO1;
assign R21C21_GB60 = R21C22_GBO1;
assign R21C22_GB60 = R21C22_GBO1;
assign R21C23_GB60 = R21C22_GBO1;
assign R21C24_GB60 = R21C22_GBO1;
assign R22C21_GB60 = R22C22_GBO1;
assign R22C22_GB60 = R22C22_GBO1;
assign R22C23_GB60 = R22C22_GBO1;
assign R22C24_GB60 = R22C22_GBO1;
assign R23C21_GB60 = R23C22_GBO1;
assign R23C22_GB60 = R23C22_GBO1;
assign R23C23_GB60 = R23C22_GBO1;
assign R23C24_GB60 = R23C22_GBO1;
assign R24C21_GB60 = R24C22_GBO1;
assign R24C22_GB60 = R24C22_GBO1;
assign R24C23_GB60 = R24C22_GBO1;
assign R24C24_GB60 = R24C22_GBO1;
assign R25C21_GB60 = R25C22_GBO1;
assign R25C22_GB60 = R25C22_GBO1;
assign R25C23_GB60 = R25C22_GBO1;
assign R25C24_GB60 = R25C22_GBO1;
assign R26C21_GB60 = R26C22_GBO1;
assign R26C22_GB60 = R26C22_GBO1;
assign R26C23_GB60 = R26C22_GBO1;
assign R26C24_GB60 = R26C22_GBO1;
assign R27C21_GB60 = R27C22_GBO1;
assign R27C22_GB60 = R27C22_GBO1;
assign R27C23_GB60 = R27C22_GBO1;
assign R27C24_GB60 = R27C22_GBO1;
assign R11C25_GB60 = R11C26_GBO1;
assign R11C26_GB60 = R11C26_GBO1;
assign R11C27_GB60 = R11C26_GBO1;
assign R11C28_GB60 = R11C26_GBO1;
assign R12C25_GB60 = R12C26_GBO1;
assign R12C26_GB60 = R12C26_GBO1;
assign R12C27_GB60 = R12C26_GBO1;
assign R12C28_GB60 = R12C26_GBO1;
assign R13C25_GB60 = R13C26_GBO1;
assign R13C26_GB60 = R13C26_GBO1;
assign R13C27_GB60 = R13C26_GBO1;
assign R13C28_GB60 = R13C26_GBO1;
assign R14C25_GB60 = R14C26_GBO1;
assign R14C26_GB60 = R14C26_GBO1;
assign R14C27_GB60 = R14C26_GBO1;
assign R14C28_GB60 = R14C26_GBO1;
assign R15C25_GB60 = R15C26_GBO1;
assign R15C26_GB60 = R15C26_GBO1;
assign R15C27_GB60 = R15C26_GBO1;
assign R15C28_GB60 = R15C26_GBO1;
assign R16C25_GB60 = R16C26_GBO1;
assign R16C26_GB60 = R16C26_GBO1;
assign R16C27_GB60 = R16C26_GBO1;
assign R16C28_GB60 = R16C26_GBO1;
assign R17C25_GB60 = R17C26_GBO1;
assign R17C26_GB60 = R17C26_GBO1;
assign R17C27_GB60 = R17C26_GBO1;
assign R17C28_GB60 = R17C26_GBO1;
assign R18C25_GB60 = R18C26_GBO1;
assign R18C26_GB60 = R18C26_GBO1;
assign R18C27_GB60 = R18C26_GBO1;
assign R18C28_GB60 = R18C26_GBO1;
assign R20C25_GB60 = R20C26_GBO1;
assign R20C26_GB60 = R20C26_GBO1;
assign R20C27_GB60 = R20C26_GBO1;
assign R20C28_GB60 = R20C26_GBO1;
assign R21C25_GB60 = R21C26_GBO1;
assign R21C26_GB60 = R21C26_GBO1;
assign R21C27_GB60 = R21C26_GBO1;
assign R21C28_GB60 = R21C26_GBO1;
assign R22C25_GB60 = R22C26_GBO1;
assign R22C26_GB60 = R22C26_GBO1;
assign R22C27_GB60 = R22C26_GBO1;
assign R22C28_GB60 = R22C26_GBO1;
assign R23C25_GB60 = R23C26_GBO1;
assign R23C26_GB60 = R23C26_GBO1;
assign R23C27_GB60 = R23C26_GBO1;
assign R23C28_GB60 = R23C26_GBO1;
assign R24C25_GB60 = R24C26_GBO1;
assign R24C26_GB60 = R24C26_GBO1;
assign R24C27_GB60 = R24C26_GBO1;
assign R24C28_GB60 = R24C26_GBO1;
assign R25C25_GB60 = R25C26_GBO1;
assign R25C26_GB60 = R25C26_GBO1;
assign R25C27_GB60 = R25C26_GBO1;
assign R25C28_GB60 = R25C26_GBO1;
assign R26C25_GB60 = R26C26_GBO1;
assign R26C26_GB60 = R26C26_GBO1;
assign R26C27_GB60 = R26C26_GBO1;
assign R26C28_GB60 = R26C26_GBO1;
assign R27C25_GB60 = R27C26_GBO1;
assign R27C26_GB60 = R27C26_GBO1;
assign R27C27_GB60 = R27C26_GBO1;
assign R27C28_GB60 = R27C26_GBO1;
assign R11C2_GB70 = R11C1_GBO1;
assign R11C3_GB70 = R11C1_GBO1;
assign R12C2_GB70 = R12C1_GBO1;
assign R12C3_GB70 = R12C1_GBO1;
assign R13C2_GB70 = R13C1_GBO1;
assign R13C3_GB70 = R13C1_GBO1;
assign R14C2_GB70 = R14C1_GBO1;
assign R14C3_GB70 = R14C1_GBO1;
assign R15C2_GB70 = R15C1_GBO1;
assign R15C3_GB70 = R15C1_GBO1;
assign R16C2_GB70 = R16C1_GBO1;
assign R16C3_GB70 = R16C1_GBO1;
assign R17C2_GB70 = R17C1_GBO1;
assign R17C3_GB70 = R17C1_GBO1;
assign R18C2_GB70 = R18C1_GBO1;
assign R18C3_GB70 = R18C1_GBO1;
assign R20C2_GB70 = R20C1_GBO1;
assign R20C3_GB70 = R20C1_GBO1;
assign R21C2_GB70 = R21C1_GBO1;
assign R21C3_GB70 = R21C1_GBO1;
assign R22C2_GB70 = R22C1_GBO1;
assign R22C3_GB70 = R22C1_GBO1;
assign R23C2_GB70 = R23C1_GBO1;
assign R23C3_GB70 = R23C1_GBO1;
assign R24C2_GB70 = R24C1_GBO1;
assign R24C3_GB70 = R24C1_GBO1;
assign R25C2_GB70 = R25C1_GBO1;
assign R25C3_GB70 = R25C1_GBO1;
assign R26C2_GB70 = R26C1_GBO1;
assign R26C3_GB70 = R26C1_GBO1;
assign R27C2_GB70 = R27C1_GBO1;
assign R27C3_GB70 = R27C1_GBO1;
assign R11C4_GB70 = R11C5_GBO1;
assign R11C5_GB70 = R11C5_GBO1;
assign R11C6_GB70 = R11C5_GBO1;
assign R11C7_GB70 = R11C5_GBO1;
assign R12C4_GB70 = R12C5_GBO1;
assign R12C5_GB70 = R12C5_GBO1;
assign R12C6_GB70 = R12C5_GBO1;
assign R12C7_GB70 = R12C5_GBO1;
assign R13C4_GB70 = R13C5_GBO1;
assign R13C5_GB70 = R13C5_GBO1;
assign R13C6_GB70 = R13C5_GBO1;
assign R13C7_GB70 = R13C5_GBO1;
assign R14C4_GB70 = R14C5_GBO1;
assign R14C5_GB70 = R14C5_GBO1;
assign R14C6_GB70 = R14C5_GBO1;
assign R14C7_GB70 = R14C5_GBO1;
assign R15C4_GB70 = R15C5_GBO1;
assign R15C5_GB70 = R15C5_GBO1;
assign R15C6_GB70 = R15C5_GBO1;
assign R15C7_GB70 = R15C5_GBO1;
assign R16C4_GB70 = R16C5_GBO1;
assign R16C5_GB70 = R16C5_GBO1;
assign R16C6_GB70 = R16C5_GBO1;
assign R16C7_GB70 = R16C5_GBO1;
assign R17C4_GB70 = R17C5_GBO1;
assign R17C5_GB70 = R17C5_GBO1;
assign R17C6_GB70 = R17C5_GBO1;
assign R17C7_GB70 = R17C5_GBO1;
assign R18C4_GB70 = R18C5_GBO1;
assign R18C5_GB70 = R18C5_GBO1;
assign R18C6_GB70 = R18C5_GBO1;
assign R18C7_GB70 = R18C5_GBO1;
assign R20C4_GB70 = R20C5_GBO1;
assign R20C5_GB70 = R20C5_GBO1;
assign R20C6_GB70 = R20C5_GBO1;
assign R20C7_GB70 = R20C5_GBO1;
assign R21C4_GB70 = R21C5_GBO1;
assign R21C5_GB70 = R21C5_GBO1;
assign R21C6_GB70 = R21C5_GBO1;
assign R21C7_GB70 = R21C5_GBO1;
assign R22C4_GB70 = R22C5_GBO1;
assign R22C5_GB70 = R22C5_GBO1;
assign R22C6_GB70 = R22C5_GBO1;
assign R22C7_GB70 = R22C5_GBO1;
assign R23C4_GB70 = R23C5_GBO1;
assign R23C5_GB70 = R23C5_GBO1;
assign R23C6_GB70 = R23C5_GBO1;
assign R23C7_GB70 = R23C5_GBO1;
assign R24C4_GB70 = R24C5_GBO1;
assign R24C5_GB70 = R24C5_GBO1;
assign R24C6_GB70 = R24C5_GBO1;
assign R24C7_GB70 = R24C5_GBO1;
assign R25C4_GB70 = R25C5_GBO1;
assign R25C5_GB70 = R25C5_GBO1;
assign R25C6_GB70 = R25C5_GBO1;
assign R25C7_GB70 = R25C5_GBO1;
assign R26C4_GB70 = R26C5_GBO1;
assign R26C5_GB70 = R26C5_GBO1;
assign R26C6_GB70 = R26C5_GBO1;
assign R26C7_GB70 = R26C5_GBO1;
assign R27C4_GB70 = R27C5_GBO1;
assign R27C5_GB70 = R27C5_GBO1;
assign R27C6_GB70 = R27C5_GBO1;
assign R27C7_GB70 = R27C5_GBO1;
assign R11C9_GB70 = R11C9_GBO1;
assign R11C10_GB70 = R11C9_GBO1;
assign R11C11_GB70 = R11C9_GBO1;
assign R11C8_GB70 = R11C9_GBO1;
assign R12C9_GB70 = R12C9_GBO1;
assign R12C10_GB70 = R12C9_GBO1;
assign R12C11_GB70 = R12C9_GBO1;
assign R12C8_GB70 = R12C9_GBO1;
assign R13C9_GB70 = R13C9_GBO1;
assign R13C10_GB70 = R13C9_GBO1;
assign R13C11_GB70 = R13C9_GBO1;
assign R13C8_GB70 = R13C9_GBO1;
assign R14C9_GB70 = R14C9_GBO1;
assign R14C10_GB70 = R14C9_GBO1;
assign R14C11_GB70 = R14C9_GBO1;
assign R14C8_GB70 = R14C9_GBO1;
assign R15C9_GB70 = R15C9_GBO1;
assign R15C10_GB70 = R15C9_GBO1;
assign R15C11_GB70 = R15C9_GBO1;
assign R15C8_GB70 = R15C9_GBO1;
assign R16C9_GB70 = R16C9_GBO1;
assign R16C10_GB70 = R16C9_GBO1;
assign R16C11_GB70 = R16C9_GBO1;
assign R16C8_GB70 = R16C9_GBO1;
assign R17C9_GB70 = R17C9_GBO1;
assign R17C10_GB70 = R17C9_GBO1;
assign R17C11_GB70 = R17C9_GBO1;
assign R17C8_GB70 = R17C9_GBO1;
assign R18C9_GB70 = R18C9_GBO1;
assign R18C10_GB70 = R18C9_GBO1;
assign R18C11_GB70 = R18C9_GBO1;
assign R18C8_GB70 = R18C9_GBO1;
assign R20C9_GB70 = R20C9_GBO1;
assign R20C10_GB70 = R20C9_GBO1;
assign R20C11_GB70 = R20C9_GBO1;
assign R20C8_GB70 = R20C9_GBO1;
assign R21C9_GB70 = R21C9_GBO1;
assign R21C10_GB70 = R21C9_GBO1;
assign R21C11_GB70 = R21C9_GBO1;
assign R21C8_GB70 = R21C9_GBO1;
assign R22C9_GB70 = R22C9_GBO1;
assign R22C10_GB70 = R22C9_GBO1;
assign R22C11_GB70 = R22C9_GBO1;
assign R22C8_GB70 = R22C9_GBO1;
assign R23C9_GB70 = R23C9_GBO1;
assign R23C10_GB70 = R23C9_GBO1;
assign R23C11_GB70 = R23C9_GBO1;
assign R23C8_GB70 = R23C9_GBO1;
assign R24C9_GB70 = R24C9_GBO1;
assign R24C10_GB70 = R24C9_GBO1;
assign R24C11_GB70 = R24C9_GBO1;
assign R24C8_GB70 = R24C9_GBO1;
assign R25C9_GB70 = R25C9_GBO1;
assign R25C10_GB70 = R25C9_GBO1;
assign R25C11_GB70 = R25C9_GBO1;
assign R25C8_GB70 = R25C9_GBO1;
assign R26C9_GB70 = R26C9_GBO1;
assign R26C10_GB70 = R26C9_GBO1;
assign R26C11_GB70 = R26C9_GBO1;
assign R26C8_GB70 = R26C9_GBO1;
assign R27C9_GB70 = R27C9_GBO1;
assign R27C10_GB70 = R27C9_GBO1;
assign R27C11_GB70 = R27C9_GBO1;
assign R27C8_GB70 = R27C9_GBO1;
assign R11C12_GB70 = R11C13_GBO1;
assign R11C13_GB70 = R11C13_GBO1;
assign R11C14_GB70 = R11C13_GBO1;
assign R11C15_GB70 = R11C13_GBO1;
assign R12C12_GB70 = R12C13_GBO1;
assign R12C13_GB70 = R12C13_GBO1;
assign R12C14_GB70 = R12C13_GBO1;
assign R12C15_GB70 = R12C13_GBO1;
assign R13C12_GB70 = R13C13_GBO1;
assign R13C13_GB70 = R13C13_GBO1;
assign R13C14_GB70 = R13C13_GBO1;
assign R13C15_GB70 = R13C13_GBO1;
assign R14C12_GB70 = R14C13_GBO1;
assign R14C13_GB70 = R14C13_GBO1;
assign R14C14_GB70 = R14C13_GBO1;
assign R14C15_GB70 = R14C13_GBO1;
assign R15C12_GB70 = R15C13_GBO1;
assign R15C13_GB70 = R15C13_GBO1;
assign R15C14_GB70 = R15C13_GBO1;
assign R15C15_GB70 = R15C13_GBO1;
assign R16C12_GB70 = R16C13_GBO1;
assign R16C13_GB70 = R16C13_GBO1;
assign R16C14_GB70 = R16C13_GBO1;
assign R16C15_GB70 = R16C13_GBO1;
assign R17C12_GB70 = R17C13_GBO1;
assign R17C13_GB70 = R17C13_GBO1;
assign R17C14_GB70 = R17C13_GBO1;
assign R17C15_GB70 = R17C13_GBO1;
assign R18C12_GB70 = R18C13_GBO1;
assign R18C13_GB70 = R18C13_GBO1;
assign R18C14_GB70 = R18C13_GBO1;
assign R18C15_GB70 = R18C13_GBO1;
assign R20C12_GB70 = R20C13_GBO1;
assign R20C13_GB70 = R20C13_GBO1;
assign R20C14_GB70 = R20C13_GBO1;
assign R20C15_GB70 = R20C13_GBO1;
assign R21C12_GB70 = R21C13_GBO1;
assign R21C13_GB70 = R21C13_GBO1;
assign R21C14_GB70 = R21C13_GBO1;
assign R21C15_GB70 = R21C13_GBO1;
assign R22C12_GB70 = R22C13_GBO1;
assign R22C13_GB70 = R22C13_GBO1;
assign R22C14_GB70 = R22C13_GBO1;
assign R22C15_GB70 = R22C13_GBO1;
assign R23C12_GB70 = R23C13_GBO1;
assign R23C13_GB70 = R23C13_GBO1;
assign R23C14_GB70 = R23C13_GBO1;
assign R23C15_GB70 = R23C13_GBO1;
assign R24C12_GB70 = R24C13_GBO1;
assign R24C13_GB70 = R24C13_GBO1;
assign R24C14_GB70 = R24C13_GBO1;
assign R24C15_GB70 = R24C13_GBO1;
assign R25C12_GB70 = R25C13_GBO1;
assign R25C13_GB70 = R25C13_GBO1;
assign R25C14_GB70 = R25C13_GBO1;
assign R25C15_GB70 = R25C13_GBO1;
assign R26C12_GB70 = R26C13_GBO1;
assign R26C13_GB70 = R26C13_GBO1;
assign R26C14_GB70 = R26C13_GBO1;
assign R26C15_GB70 = R26C13_GBO1;
assign R27C12_GB70 = R27C13_GBO1;
assign R27C13_GB70 = R27C13_GBO1;
assign R27C14_GB70 = R27C13_GBO1;
assign R27C15_GB70 = R27C13_GBO1;
assign R11C17_GB70 = R11C17_GBO1;
assign R11C18_GB70 = R11C17_GBO1;
assign R11C19_GB70 = R11C17_GBO1;
assign R11C16_GB70 = R11C17_GBO1;
assign R12C17_GB70 = R12C17_GBO1;
assign R12C18_GB70 = R12C17_GBO1;
assign R12C19_GB70 = R12C17_GBO1;
assign R12C16_GB70 = R12C17_GBO1;
assign R13C17_GB70 = R13C17_GBO1;
assign R13C18_GB70 = R13C17_GBO1;
assign R13C19_GB70 = R13C17_GBO1;
assign R13C16_GB70 = R13C17_GBO1;
assign R14C17_GB70 = R14C17_GBO1;
assign R14C18_GB70 = R14C17_GBO1;
assign R14C19_GB70 = R14C17_GBO1;
assign R14C16_GB70 = R14C17_GBO1;
assign R15C17_GB70 = R15C17_GBO1;
assign R15C18_GB70 = R15C17_GBO1;
assign R15C19_GB70 = R15C17_GBO1;
assign R15C16_GB70 = R15C17_GBO1;
assign R16C17_GB70 = R16C17_GBO1;
assign R16C18_GB70 = R16C17_GBO1;
assign R16C19_GB70 = R16C17_GBO1;
assign R16C16_GB70 = R16C17_GBO1;
assign R17C17_GB70 = R17C17_GBO1;
assign R17C18_GB70 = R17C17_GBO1;
assign R17C19_GB70 = R17C17_GBO1;
assign R17C16_GB70 = R17C17_GBO1;
assign R18C17_GB70 = R18C17_GBO1;
assign R18C18_GB70 = R18C17_GBO1;
assign R18C19_GB70 = R18C17_GBO1;
assign R18C16_GB70 = R18C17_GBO1;
assign R20C17_GB70 = R20C17_GBO1;
assign R20C18_GB70 = R20C17_GBO1;
assign R20C19_GB70 = R20C17_GBO1;
assign R20C16_GB70 = R20C17_GBO1;
assign R21C17_GB70 = R21C17_GBO1;
assign R21C18_GB70 = R21C17_GBO1;
assign R21C19_GB70 = R21C17_GBO1;
assign R21C16_GB70 = R21C17_GBO1;
assign R22C17_GB70 = R22C17_GBO1;
assign R22C18_GB70 = R22C17_GBO1;
assign R22C19_GB70 = R22C17_GBO1;
assign R22C16_GB70 = R22C17_GBO1;
assign R23C17_GB70 = R23C17_GBO1;
assign R23C18_GB70 = R23C17_GBO1;
assign R23C19_GB70 = R23C17_GBO1;
assign R23C16_GB70 = R23C17_GBO1;
assign R24C17_GB70 = R24C17_GBO1;
assign R24C18_GB70 = R24C17_GBO1;
assign R24C19_GB70 = R24C17_GBO1;
assign R24C16_GB70 = R24C17_GBO1;
assign R25C17_GB70 = R25C17_GBO1;
assign R25C18_GB70 = R25C17_GBO1;
assign R25C19_GB70 = R25C17_GBO1;
assign R25C16_GB70 = R25C17_GBO1;
assign R26C17_GB70 = R26C17_GBO1;
assign R26C18_GB70 = R26C17_GBO1;
assign R26C19_GB70 = R26C17_GBO1;
assign R26C16_GB70 = R26C17_GBO1;
assign R27C17_GB70 = R27C17_GBO1;
assign R27C18_GB70 = R27C17_GBO1;
assign R27C19_GB70 = R27C17_GBO1;
assign R27C16_GB70 = R27C17_GBO1;
assign R11C20_GB70 = R11C21_GBO1;
assign R11C21_GB70 = R11C21_GBO1;
assign R11C22_GB70 = R11C21_GBO1;
assign R11C23_GB70 = R11C21_GBO1;
assign R12C20_GB70 = R12C21_GBO1;
assign R12C21_GB70 = R12C21_GBO1;
assign R12C22_GB70 = R12C21_GBO1;
assign R12C23_GB70 = R12C21_GBO1;
assign R13C20_GB70 = R13C21_GBO1;
assign R13C21_GB70 = R13C21_GBO1;
assign R13C22_GB70 = R13C21_GBO1;
assign R13C23_GB70 = R13C21_GBO1;
assign R14C20_GB70 = R14C21_GBO1;
assign R14C21_GB70 = R14C21_GBO1;
assign R14C22_GB70 = R14C21_GBO1;
assign R14C23_GB70 = R14C21_GBO1;
assign R15C20_GB70 = R15C21_GBO1;
assign R15C21_GB70 = R15C21_GBO1;
assign R15C22_GB70 = R15C21_GBO1;
assign R15C23_GB70 = R15C21_GBO1;
assign R16C20_GB70 = R16C21_GBO1;
assign R16C21_GB70 = R16C21_GBO1;
assign R16C22_GB70 = R16C21_GBO1;
assign R16C23_GB70 = R16C21_GBO1;
assign R17C20_GB70 = R17C21_GBO1;
assign R17C21_GB70 = R17C21_GBO1;
assign R17C22_GB70 = R17C21_GBO1;
assign R17C23_GB70 = R17C21_GBO1;
assign R18C20_GB70 = R18C21_GBO1;
assign R18C21_GB70 = R18C21_GBO1;
assign R18C22_GB70 = R18C21_GBO1;
assign R18C23_GB70 = R18C21_GBO1;
assign R20C20_GB70 = R20C21_GBO1;
assign R20C21_GB70 = R20C21_GBO1;
assign R20C22_GB70 = R20C21_GBO1;
assign R20C23_GB70 = R20C21_GBO1;
assign R21C20_GB70 = R21C21_GBO1;
assign R21C21_GB70 = R21C21_GBO1;
assign R21C22_GB70 = R21C21_GBO1;
assign R21C23_GB70 = R21C21_GBO1;
assign R22C20_GB70 = R22C21_GBO1;
assign R22C21_GB70 = R22C21_GBO1;
assign R22C22_GB70 = R22C21_GBO1;
assign R22C23_GB70 = R22C21_GBO1;
assign R23C20_GB70 = R23C21_GBO1;
assign R23C21_GB70 = R23C21_GBO1;
assign R23C22_GB70 = R23C21_GBO1;
assign R23C23_GB70 = R23C21_GBO1;
assign R24C20_GB70 = R24C21_GBO1;
assign R24C21_GB70 = R24C21_GBO1;
assign R24C22_GB70 = R24C21_GBO1;
assign R24C23_GB70 = R24C21_GBO1;
assign R25C20_GB70 = R25C21_GBO1;
assign R25C21_GB70 = R25C21_GBO1;
assign R25C22_GB70 = R25C21_GBO1;
assign R25C23_GB70 = R25C21_GBO1;
assign R26C20_GB70 = R26C21_GBO1;
assign R26C21_GB70 = R26C21_GBO1;
assign R26C22_GB70 = R26C21_GBO1;
assign R26C23_GB70 = R26C21_GBO1;
assign R27C20_GB70 = R27C21_GBO1;
assign R27C21_GB70 = R27C21_GBO1;
assign R27C22_GB70 = R27C21_GBO1;
assign R27C23_GB70 = R27C21_GBO1;
assign R11C24_GB70 = R11C25_GBO1;
assign R11C25_GB70 = R11C25_GBO1;
assign R11C26_GB70 = R11C25_GBO1;
assign R11C27_GB70 = R11C25_GBO1;
assign R11C28_GB70 = R11C25_GBO1;
assign R12C24_GB70 = R12C25_GBO1;
assign R12C25_GB70 = R12C25_GBO1;
assign R12C26_GB70 = R12C25_GBO1;
assign R12C27_GB70 = R12C25_GBO1;
assign R12C28_GB70 = R12C25_GBO1;
assign R13C24_GB70 = R13C25_GBO1;
assign R13C25_GB70 = R13C25_GBO1;
assign R13C26_GB70 = R13C25_GBO1;
assign R13C27_GB70 = R13C25_GBO1;
assign R13C28_GB70 = R13C25_GBO1;
assign R14C24_GB70 = R14C25_GBO1;
assign R14C25_GB70 = R14C25_GBO1;
assign R14C26_GB70 = R14C25_GBO1;
assign R14C27_GB70 = R14C25_GBO1;
assign R14C28_GB70 = R14C25_GBO1;
assign R15C24_GB70 = R15C25_GBO1;
assign R15C25_GB70 = R15C25_GBO1;
assign R15C26_GB70 = R15C25_GBO1;
assign R15C27_GB70 = R15C25_GBO1;
assign R15C28_GB70 = R15C25_GBO1;
assign R16C24_GB70 = R16C25_GBO1;
assign R16C25_GB70 = R16C25_GBO1;
assign R16C26_GB70 = R16C25_GBO1;
assign R16C27_GB70 = R16C25_GBO1;
assign R16C28_GB70 = R16C25_GBO1;
assign R17C24_GB70 = R17C25_GBO1;
assign R17C25_GB70 = R17C25_GBO1;
assign R17C26_GB70 = R17C25_GBO1;
assign R17C27_GB70 = R17C25_GBO1;
assign R17C28_GB70 = R17C25_GBO1;
assign R18C24_GB70 = R18C25_GBO1;
assign R18C25_GB70 = R18C25_GBO1;
assign R18C26_GB70 = R18C25_GBO1;
assign R18C27_GB70 = R18C25_GBO1;
assign R18C28_GB70 = R18C25_GBO1;
assign R20C24_GB70 = R20C25_GBO1;
assign R20C25_GB70 = R20C25_GBO1;
assign R20C26_GB70 = R20C25_GBO1;
assign R20C27_GB70 = R20C25_GBO1;
assign R20C28_GB70 = R20C25_GBO1;
assign R21C24_GB70 = R21C25_GBO1;
assign R21C25_GB70 = R21C25_GBO1;
assign R21C26_GB70 = R21C25_GBO1;
assign R21C27_GB70 = R21C25_GBO1;
assign R21C28_GB70 = R21C25_GBO1;
assign R22C24_GB70 = R22C25_GBO1;
assign R22C25_GB70 = R22C25_GBO1;
assign R22C26_GB70 = R22C25_GBO1;
assign R22C27_GB70 = R22C25_GBO1;
assign R22C28_GB70 = R22C25_GBO1;
assign R23C24_GB70 = R23C25_GBO1;
assign R23C25_GB70 = R23C25_GBO1;
assign R23C26_GB70 = R23C25_GBO1;
assign R23C27_GB70 = R23C25_GBO1;
assign R23C28_GB70 = R23C25_GBO1;
assign R24C24_GB70 = R24C25_GBO1;
assign R24C25_GB70 = R24C25_GBO1;
assign R24C26_GB70 = R24C25_GBO1;
assign R24C27_GB70 = R24C25_GBO1;
assign R24C28_GB70 = R24C25_GBO1;
assign R25C24_GB70 = R25C25_GBO1;
assign R25C25_GB70 = R25C25_GBO1;
assign R25C26_GB70 = R25C25_GBO1;
assign R25C27_GB70 = R25C25_GBO1;
assign R25C28_GB70 = R25C25_GBO1;
assign R26C24_GB70 = R26C25_GBO1;
assign R26C25_GB70 = R26C25_GBO1;
assign R26C26_GB70 = R26C25_GBO1;
assign R26C27_GB70 = R26C25_GBO1;
assign R26C28_GB70 = R26C25_GBO1;
assign R27C24_GB70 = R27C25_GBO1;
assign R27C25_GB70 = R27C25_GBO1;
assign R27C26_GB70 = R27C25_GBO1;
assign R27C27_GB70 = R27C25_GBO1;
assign R27C28_GB70 = R27C25_GBO1;
assign R2C33_GB00 = R2C32_GBO0;
assign R2C34_GB00 = R2C32_GBO0;
assign R2C29_GB00 = R2C32_GBO0;
assign R2C30_GB00 = R2C32_GBO0;
assign R2C31_GB00 = R2C32_GBO0;
assign R2C32_GB00 = R2C32_GBO0;
assign R3C33_GB00 = R3C32_GBO0;
assign R3C34_GB00 = R3C32_GBO0;
assign R3C29_GB00 = R3C32_GBO0;
assign R3C30_GB00 = R3C32_GBO0;
assign R3C31_GB00 = R3C32_GBO0;
assign R3C32_GB00 = R3C32_GBO0;
assign R4C33_GB00 = R4C32_GBO0;
assign R4C34_GB00 = R4C32_GBO0;
assign R4C29_GB00 = R4C32_GBO0;
assign R4C30_GB00 = R4C32_GBO0;
assign R4C31_GB00 = R4C32_GBO0;
assign R4C32_GB00 = R4C32_GBO0;
assign R5C33_GB00 = R5C32_GBO0;
assign R5C34_GB00 = R5C32_GBO0;
assign R5C29_GB00 = R5C32_GBO0;
assign R5C30_GB00 = R5C32_GBO0;
assign R5C31_GB00 = R5C32_GBO0;
assign R5C32_GB00 = R5C32_GBO0;
assign R6C33_GB00 = R6C32_GBO0;
assign R6C34_GB00 = R6C32_GBO0;
assign R6C29_GB00 = R6C32_GBO0;
assign R6C30_GB00 = R6C32_GBO0;
assign R6C31_GB00 = R6C32_GBO0;
assign R6C32_GB00 = R6C32_GBO0;
assign R7C33_GB00 = R7C32_GBO0;
assign R7C34_GB00 = R7C32_GBO0;
assign R7C29_GB00 = R7C32_GBO0;
assign R7C30_GB00 = R7C32_GBO0;
assign R7C31_GB00 = R7C32_GBO0;
assign R7C32_GB00 = R7C32_GBO0;
assign R8C33_GB00 = R8C32_GBO0;
assign R8C34_GB00 = R8C32_GBO0;
assign R8C29_GB00 = R8C32_GBO0;
assign R8C30_GB00 = R8C32_GBO0;
assign R8C31_GB00 = R8C32_GBO0;
assign R8C32_GB00 = R8C32_GBO0;
assign R9C33_GB00 = R9C32_GBO0;
assign R9C34_GB00 = R9C32_GBO0;
assign R9C29_GB00 = R9C32_GBO0;
assign R9C30_GB00 = R9C32_GBO0;
assign R9C31_GB00 = R9C32_GBO0;
assign R9C32_GB00 = R9C32_GBO0;
assign R2C35_GB00 = R2C36_GBO0;
assign R2C36_GB00 = R2C36_GBO0;
assign R2C37_GB00 = R2C36_GBO0;
assign R2C38_GB00 = R2C36_GBO0;
assign R3C35_GB00 = R3C36_GBO0;
assign R3C36_GB00 = R3C36_GBO0;
assign R3C37_GB00 = R3C36_GBO0;
assign R3C38_GB00 = R3C36_GBO0;
assign R4C35_GB00 = R4C36_GBO0;
assign R4C36_GB00 = R4C36_GBO0;
assign R4C37_GB00 = R4C36_GBO0;
assign R4C38_GB00 = R4C36_GBO0;
assign R5C35_GB00 = R5C36_GBO0;
assign R5C36_GB00 = R5C36_GBO0;
assign R5C37_GB00 = R5C36_GBO0;
assign R5C38_GB00 = R5C36_GBO0;
assign R6C35_GB00 = R6C36_GBO0;
assign R6C36_GB00 = R6C36_GBO0;
assign R6C37_GB00 = R6C36_GBO0;
assign R6C38_GB00 = R6C36_GBO0;
assign R7C35_GB00 = R7C36_GBO0;
assign R7C36_GB00 = R7C36_GBO0;
assign R7C37_GB00 = R7C36_GBO0;
assign R7C38_GB00 = R7C36_GBO0;
assign R8C35_GB00 = R8C36_GBO0;
assign R8C36_GB00 = R8C36_GBO0;
assign R8C37_GB00 = R8C36_GBO0;
assign R8C38_GB00 = R8C36_GBO0;
assign R9C35_GB00 = R9C36_GBO0;
assign R9C36_GB00 = R9C36_GBO0;
assign R9C37_GB00 = R9C36_GBO0;
assign R9C38_GB00 = R9C36_GBO0;
assign R2C41_GB00 = R2C40_GBO0;
assign R2C42_GB00 = R2C40_GBO0;
assign R2C39_GB00 = R2C40_GBO0;
assign R2C40_GB00 = R2C40_GBO0;
assign R3C41_GB00 = R3C40_GBO0;
assign R3C42_GB00 = R3C40_GBO0;
assign R3C39_GB00 = R3C40_GBO0;
assign R3C40_GB00 = R3C40_GBO0;
assign R4C41_GB00 = R4C40_GBO0;
assign R4C42_GB00 = R4C40_GBO0;
assign R4C39_GB00 = R4C40_GBO0;
assign R4C40_GB00 = R4C40_GBO0;
assign R5C41_GB00 = R5C40_GBO0;
assign R5C42_GB00 = R5C40_GBO0;
assign R5C39_GB00 = R5C40_GBO0;
assign R5C40_GB00 = R5C40_GBO0;
assign R6C41_GB00 = R6C40_GBO0;
assign R6C42_GB00 = R6C40_GBO0;
assign R6C39_GB00 = R6C40_GBO0;
assign R6C40_GB00 = R6C40_GBO0;
assign R7C41_GB00 = R7C40_GBO0;
assign R7C42_GB00 = R7C40_GBO0;
assign R7C39_GB00 = R7C40_GBO0;
assign R7C40_GB00 = R7C40_GBO0;
assign R8C41_GB00 = R8C40_GBO0;
assign R8C42_GB00 = R8C40_GBO0;
assign R8C39_GB00 = R8C40_GBO0;
assign R8C40_GB00 = R8C40_GBO0;
assign R9C41_GB00 = R9C40_GBO0;
assign R9C42_GB00 = R9C40_GBO0;
assign R9C39_GB00 = R9C40_GBO0;
assign R9C40_GB00 = R9C40_GBO0;
assign R2C43_GB00 = R2C44_GBO0;
assign R2C44_GB00 = R2C44_GBO0;
assign R2C45_GB00 = R2C44_GBO0;
assign R2C46_GB00 = R2C44_GBO0;
assign R3C43_GB00 = R3C44_GBO0;
assign R3C44_GB00 = R3C44_GBO0;
assign R3C45_GB00 = R3C44_GBO0;
assign R3C46_GB00 = R3C44_GBO0;
assign R4C43_GB00 = R4C44_GBO0;
assign R4C44_GB00 = R4C44_GBO0;
assign R4C45_GB00 = R4C44_GBO0;
assign R4C46_GB00 = R4C44_GBO0;
assign R5C43_GB00 = R5C44_GBO0;
assign R5C44_GB00 = R5C44_GBO0;
assign R5C45_GB00 = R5C44_GBO0;
assign R5C46_GB00 = R5C44_GBO0;
assign R6C43_GB00 = R6C44_GBO0;
assign R6C44_GB00 = R6C44_GBO0;
assign R6C45_GB00 = R6C44_GBO0;
assign R6C46_GB00 = R6C44_GBO0;
assign R7C43_GB00 = R7C44_GBO0;
assign R7C44_GB00 = R7C44_GBO0;
assign R7C45_GB00 = R7C44_GBO0;
assign R7C46_GB00 = R7C44_GBO0;
assign R8C43_GB00 = R8C44_GBO0;
assign R8C44_GB00 = R8C44_GBO0;
assign R8C45_GB00 = R8C44_GBO0;
assign R8C46_GB00 = R8C44_GBO0;
assign R9C43_GB00 = R9C44_GBO0;
assign R9C44_GB00 = R9C44_GBO0;
assign R9C45_GB00 = R9C44_GBO0;
assign R9C46_GB00 = R9C44_GBO0;
assign R2C33_GB10 = R2C31_GBO0;
assign R2C29_GB10 = R2C31_GBO0;
assign R2C30_GB10 = R2C31_GBO0;
assign R2C31_GB10 = R2C31_GBO0;
assign R2C32_GB10 = R2C31_GBO0;
assign R3C33_GB10 = R3C31_GBO0;
assign R3C29_GB10 = R3C31_GBO0;
assign R3C30_GB10 = R3C31_GBO0;
assign R3C31_GB10 = R3C31_GBO0;
assign R3C32_GB10 = R3C31_GBO0;
assign R4C33_GB10 = R4C31_GBO0;
assign R4C29_GB10 = R4C31_GBO0;
assign R4C30_GB10 = R4C31_GBO0;
assign R4C31_GB10 = R4C31_GBO0;
assign R4C32_GB10 = R4C31_GBO0;
assign R5C33_GB10 = R5C31_GBO0;
assign R5C29_GB10 = R5C31_GBO0;
assign R5C30_GB10 = R5C31_GBO0;
assign R5C31_GB10 = R5C31_GBO0;
assign R5C32_GB10 = R5C31_GBO0;
assign R6C33_GB10 = R6C31_GBO0;
assign R6C29_GB10 = R6C31_GBO0;
assign R6C30_GB10 = R6C31_GBO0;
assign R6C31_GB10 = R6C31_GBO0;
assign R6C32_GB10 = R6C31_GBO0;
assign R7C33_GB10 = R7C31_GBO0;
assign R7C29_GB10 = R7C31_GBO0;
assign R7C30_GB10 = R7C31_GBO0;
assign R7C31_GB10 = R7C31_GBO0;
assign R7C32_GB10 = R7C31_GBO0;
assign R8C33_GB10 = R8C31_GBO0;
assign R8C29_GB10 = R8C31_GBO0;
assign R8C30_GB10 = R8C31_GBO0;
assign R8C31_GB10 = R8C31_GBO0;
assign R8C32_GB10 = R8C31_GBO0;
assign R9C33_GB10 = R9C31_GBO0;
assign R9C29_GB10 = R9C31_GBO0;
assign R9C30_GB10 = R9C31_GBO0;
assign R9C31_GB10 = R9C31_GBO0;
assign R9C32_GB10 = R9C31_GBO0;
assign R2C34_GB10 = R2C35_GBO0;
assign R2C35_GB10 = R2C35_GBO0;
assign R2C36_GB10 = R2C35_GBO0;
assign R2C37_GB10 = R2C35_GBO0;
assign R3C34_GB10 = R3C35_GBO0;
assign R3C35_GB10 = R3C35_GBO0;
assign R3C36_GB10 = R3C35_GBO0;
assign R3C37_GB10 = R3C35_GBO0;
assign R4C34_GB10 = R4C35_GBO0;
assign R4C35_GB10 = R4C35_GBO0;
assign R4C36_GB10 = R4C35_GBO0;
assign R4C37_GB10 = R4C35_GBO0;
assign R5C34_GB10 = R5C35_GBO0;
assign R5C35_GB10 = R5C35_GBO0;
assign R5C36_GB10 = R5C35_GBO0;
assign R5C37_GB10 = R5C35_GBO0;
assign R6C34_GB10 = R6C35_GBO0;
assign R6C35_GB10 = R6C35_GBO0;
assign R6C36_GB10 = R6C35_GBO0;
assign R6C37_GB10 = R6C35_GBO0;
assign R7C34_GB10 = R7C35_GBO0;
assign R7C35_GB10 = R7C35_GBO0;
assign R7C36_GB10 = R7C35_GBO0;
assign R7C37_GB10 = R7C35_GBO0;
assign R8C34_GB10 = R8C35_GBO0;
assign R8C35_GB10 = R8C35_GBO0;
assign R8C36_GB10 = R8C35_GBO0;
assign R8C37_GB10 = R8C35_GBO0;
assign R9C34_GB10 = R9C35_GBO0;
assign R9C35_GB10 = R9C35_GBO0;
assign R9C36_GB10 = R9C35_GBO0;
assign R9C37_GB10 = R9C35_GBO0;
assign R2C41_GB10 = R2C39_GBO0;
assign R2C38_GB10 = R2C39_GBO0;
assign R2C39_GB10 = R2C39_GBO0;
assign R2C40_GB10 = R2C39_GBO0;
assign R3C41_GB10 = R3C39_GBO0;
assign R3C38_GB10 = R3C39_GBO0;
assign R3C39_GB10 = R3C39_GBO0;
assign R3C40_GB10 = R3C39_GBO0;
assign R4C41_GB10 = R4C39_GBO0;
assign R4C38_GB10 = R4C39_GBO0;
assign R4C39_GB10 = R4C39_GBO0;
assign R4C40_GB10 = R4C39_GBO0;
assign R5C41_GB10 = R5C39_GBO0;
assign R5C38_GB10 = R5C39_GBO0;
assign R5C39_GB10 = R5C39_GBO0;
assign R5C40_GB10 = R5C39_GBO0;
assign R6C41_GB10 = R6C39_GBO0;
assign R6C38_GB10 = R6C39_GBO0;
assign R6C39_GB10 = R6C39_GBO0;
assign R6C40_GB10 = R6C39_GBO0;
assign R7C41_GB10 = R7C39_GBO0;
assign R7C38_GB10 = R7C39_GBO0;
assign R7C39_GB10 = R7C39_GBO0;
assign R7C40_GB10 = R7C39_GBO0;
assign R8C41_GB10 = R8C39_GBO0;
assign R8C38_GB10 = R8C39_GBO0;
assign R8C39_GB10 = R8C39_GBO0;
assign R8C40_GB10 = R8C39_GBO0;
assign R9C41_GB10 = R9C39_GBO0;
assign R9C38_GB10 = R9C39_GBO0;
assign R9C39_GB10 = R9C39_GBO0;
assign R9C40_GB10 = R9C39_GBO0;
assign R2C42_GB10 = R2C43_GBO0;
assign R2C43_GB10 = R2C43_GBO0;
assign R2C44_GB10 = R2C43_GBO0;
assign R2C45_GB10 = R2C43_GBO0;
assign R2C46_GB10 = R2C43_GBO0;
assign R3C42_GB10 = R3C43_GBO0;
assign R3C43_GB10 = R3C43_GBO0;
assign R3C44_GB10 = R3C43_GBO0;
assign R3C45_GB10 = R3C43_GBO0;
assign R3C46_GB10 = R3C43_GBO0;
assign R4C42_GB10 = R4C43_GBO0;
assign R4C43_GB10 = R4C43_GBO0;
assign R4C44_GB10 = R4C43_GBO0;
assign R4C45_GB10 = R4C43_GBO0;
assign R4C46_GB10 = R4C43_GBO0;
assign R5C42_GB10 = R5C43_GBO0;
assign R5C43_GB10 = R5C43_GBO0;
assign R5C44_GB10 = R5C43_GBO0;
assign R5C45_GB10 = R5C43_GBO0;
assign R5C46_GB10 = R5C43_GBO0;
assign R6C42_GB10 = R6C43_GBO0;
assign R6C43_GB10 = R6C43_GBO0;
assign R6C44_GB10 = R6C43_GBO0;
assign R6C45_GB10 = R6C43_GBO0;
assign R6C46_GB10 = R6C43_GBO0;
assign R7C42_GB10 = R7C43_GBO0;
assign R7C43_GB10 = R7C43_GBO0;
assign R7C44_GB10 = R7C43_GBO0;
assign R7C45_GB10 = R7C43_GBO0;
assign R7C46_GB10 = R7C43_GBO0;
assign R8C42_GB10 = R8C43_GBO0;
assign R8C43_GB10 = R8C43_GBO0;
assign R8C44_GB10 = R8C43_GBO0;
assign R8C45_GB10 = R8C43_GBO0;
assign R8C46_GB10 = R8C43_GBO0;
assign R9C42_GB10 = R9C43_GBO0;
assign R9C43_GB10 = R9C43_GBO0;
assign R9C44_GB10 = R9C43_GBO0;
assign R9C45_GB10 = R9C43_GBO0;
assign R9C46_GB10 = R9C43_GBO0;
assign R2C29_GB20 = R2C30_GBO0;
assign R2C30_GB20 = R2C30_GBO0;
assign R2C31_GB20 = R2C30_GBO0;
assign R2C32_GB20 = R2C30_GBO0;
assign R3C29_GB20 = R3C30_GBO0;
assign R3C30_GB20 = R3C30_GBO0;
assign R3C31_GB20 = R3C30_GBO0;
assign R3C32_GB20 = R3C30_GBO0;
assign R4C29_GB20 = R4C30_GBO0;
assign R4C30_GB20 = R4C30_GBO0;
assign R4C31_GB20 = R4C30_GBO0;
assign R4C32_GB20 = R4C30_GBO0;
assign R5C29_GB20 = R5C30_GBO0;
assign R5C30_GB20 = R5C30_GBO0;
assign R5C31_GB20 = R5C30_GBO0;
assign R5C32_GB20 = R5C30_GBO0;
assign R6C29_GB20 = R6C30_GBO0;
assign R6C30_GB20 = R6C30_GBO0;
assign R6C31_GB20 = R6C30_GBO0;
assign R6C32_GB20 = R6C30_GBO0;
assign R7C29_GB20 = R7C30_GBO0;
assign R7C30_GB20 = R7C30_GBO0;
assign R7C31_GB20 = R7C30_GBO0;
assign R7C32_GB20 = R7C30_GBO0;
assign R8C29_GB20 = R8C30_GBO0;
assign R8C30_GB20 = R8C30_GBO0;
assign R8C31_GB20 = R8C30_GBO0;
assign R8C32_GB20 = R8C30_GBO0;
assign R9C29_GB20 = R9C30_GBO0;
assign R9C30_GB20 = R9C30_GBO0;
assign R9C31_GB20 = R9C30_GBO0;
assign R9C32_GB20 = R9C30_GBO0;
assign R2C33_GB20 = R2C34_GBO0;
assign R2C34_GB20 = R2C34_GBO0;
assign R2C35_GB20 = R2C34_GBO0;
assign R2C36_GB20 = R2C34_GBO0;
assign R3C33_GB20 = R3C34_GBO0;
assign R3C34_GB20 = R3C34_GBO0;
assign R3C35_GB20 = R3C34_GBO0;
assign R3C36_GB20 = R3C34_GBO0;
assign R4C33_GB20 = R4C34_GBO0;
assign R4C34_GB20 = R4C34_GBO0;
assign R4C35_GB20 = R4C34_GBO0;
assign R4C36_GB20 = R4C34_GBO0;
assign R5C33_GB20 = R5C34_GBO0;
assign R5C34_GB20 = R5C34_GBO0;
assign R5C35_GB20 = R5C34_GBO0;
assign R5C36_GB20 = R5C34_GBO0;
assign R6C33_GB20 = R6C34_GBO0;
assign R6C34_GB20 = R6C34_GBO0;
assign R6C35_GB20 = R6C34_GBO0;
assign R6C36_GB20 = R6C34_GBO0;
assign R7C33_GB20 = R7C34_GBO0;
assign R7C34_GB20 = R7C34_GBO0;
assign R7C35_GB20 = R7C34_GBO0;
assign R7C36_GB20 = R7C34_GBO0;
assign R8C33_GB20 = R8C34_GBO0;
assign R8C34_GB20 = R8C34_GBO0;
assign R8C35_GB20 = R8C34_GBO0;
assign R8C36_GB20 = R8C34_GBO0;
assign R9C33_GB20 = R9C34_GBO0;
assign R9C34_GB20 = R9C34_GBO0;
assign R9C35_GB20 = R9C34_GBO0;
assign R9C36_GB20 = R9C34_GBO0;
assign R2C37_GB20 = R2C38_GBO0;
assign R2C38_GB20 = R2C38_GBO0;
assign R2C39_GB20 = R2C38_GBO0;
assign R2C40_GB20 = R2C38_GBO0;
assign R3C37_GB20 = R3C38_GBO0;
assign R3C38_GB20 = R3C38_GBO0;
assign R3C39_GB20 = R3C38_GBO0;
assign R3C40_GB20 = R3C38_GBO0;
assign R4C37_GB20 = R4C38_GBO0;
assign R4C38_GB20 = R4C38_GBO0;
assign R4C39_GB20 = R4C38_GBO0;
assign R4C40_GB20 = R4C38_GBO0;
assign R5C37_GB20 = R5C38_GBO0;
assign R5C38_GB20 = R5C38_GBO0;
assign R5C39_GB20 = R5C38_GBO0;
assign R5C40_GB20 = R5C38_GBO0;
assign R6C37_GB20 = R6C38_GBO0;
assign R6C38_GB20 = R6C38_GBO0;
assign R6C39_GB20 = R6C38_GBO0;
assign R6C40_GB20 = R6C38_GBO0;
assign R7C37_GB20 = R7C38_GBO0;
assign R7C38_GB20 = R7C38_GBO0;
assign R7C39_GB20 = R7C38_GBO0;
assign R7C40_GB20 = R7C38_GBO0;
assign R8C37_GB20 = R8C38_GBO0;
assign R8C38_GB20 = R8C38_GBO0;
assign R8C39_GB20 = R8C38_GBO0;
assign R8C40_GB20 = R8C38_GBO0;
assign R9C37_GB20 = R9C38_GBO0;
assign R9C38_GB20 = R9C38_GBO0;
assign R9C39_GB20 = R9C38_GBO0;
assign R9C40_GB20 = R9C38_GBO0;
assign R2C41_GB20 = R2C42_GBO0;
assign R2C42_GB20 = R2C42_GBO0;
assign R2C43_GB20 = R2C42_GBO0;
assign R2C44_GB20 = R2C42_GBO0;
assign R3C41_GB20 = R3C42_GBO0;
assign R3C42_GB20 = R3C42_GBO0;
assign R3C43_GB20 = R3C42_GBO0;
assign R3C44_GB20 = R3C42_GBO0;
assign R4C41_GB20 = R4C42_GBO0;
assign R4C42_GB20 = R4C42_GBO0;
assign R4C43_GB20 = R4C42_GBO0;
assign R4C44_GB20 = R4C42_GBO0;
assign R5C41_GB20 = R5C42_GBO0;
assign R5C42_GB20 = R5C42_GBO0;
assign R5C43_GB20 = R5C42_GBO0;
assign R5C44_GB20 = R5C42_GBO0;
assign R6C41_GB20 = R6C42_GBO0;
assign R6C42_GB20 = R6C42_GBO0;
assign R6C43_GB20 = R6C42_GBO0;
assign R6C44_GB20 = R6C42_GBO0;
assign R7C41_GB20 = R7C42_GBO0;
assign R7C42_GB20 = R7C42_GBO0;
assign R7C43_GB20 = R7C42_GBO0;
assign R7C44_GB20 = R7C42_GBO0;
assign R8C41_GB20 = R8C42_GBO0;
assign R8C42_GB20 = R8C42_GBO0;
assign R8C43_GB20 = R8C42_GBO0;
assign R8C44_GB20 = R8C42_GBO0;
assign R9C41_GB20 = R9C42_GBO0;
assign R9C42_GB20 = R9C42_GBO0;
assign R9C43_GB20 = R9C42_GBO0;
assign R9C44_GB20 = R9C42_GBO0;
assign R2C45_GB20 = R2C46_GBO0;
assign R2C46_GB20 = R2C46_GBO0;
assign R3C45_GB20 = R3C46_GBO0;
assign R3C46_GB20 = R3C46_GBO0;
assign R4C45_GB20 = R4C46_GBO0;
assign R4C46_GB20 = R4C46_GBO0;
assign R5C45_GB20 = R5C46_GBO0;
assign R5C46_GB20 = R5C46_GBO0;
assign R6C45_GB20 = R6C46_GBO0;
assign R6C46_GB20 = R6C46_GBO0;
assign R7C45_GB20 = R7C46_GBO0;
assign R7C46_GB20 = R7C46_GBO0;
assign R8C45_GB20 = R8C46_GBO0;
assign R8C46_GB20 = R8C46_GBO0;
assign R9C45_GB20 = R9C46_GBO0;
assign R9C46_GB20 = R9C46_GBO0;
assign R2C29_GB30 = R2C29_GBO0;
assign R2C30_GB30 = R2C29_GBO0;
assign R2C31_GB30 = R2C29_GBO0;
assign R3C29_GB30 = R3C29_GBO0;
assign R3C30_GB30 = R3C29_GBO0;
assign R3C31_GB30 = R3C29_GBO0;
assign R4C29_GB30 = R4C29_GBO0;
assign R4C30_GB30 = R4C29_GBO0;
assign R4C31_GB30 = R4C29_GBO0;
assign R5C29_GB30 = R5C29_GBO0;
assign R5C30_GB30 = R5C29_GBO0;
assign R5C31_GB30 = R5C29_GBO0;
assign R6C29_GB30 = R6C29_GBO0;
assign R6C30_GB30 = R6C29_GBO0;
assign R6C31_GB30 = R6C29_GBO0;
assign R7C29_GB30 = R7C29_GBO0;
assign R7C30_GB30 = R7C29_GBO0;
assign R7C31_GB30 = R7C29_GBO0;
assign R8C29_GB30 = R8C29_GBO0;
assign R8C30_GB30 = R8C29_GBO0;
assign R8C31_GB30 = R8C29_GBO0;
assign R9C29_GB30 = R9C29_GBO0;
assign R9C30_GB30 = R9C29_GBO0;
assign R9C31_GB30 = R9C29_GBO0;
assign R2C33_GB30 = R2C33_GBO0;
assign R2C34_GB30 = R2C33_GBO0;
assign R2C35_GB30 = R2C33_GBO0;
assign R2C32_GB30 = R2C33_GBO0;
assign R3C33_GB30 = R3C33_GBO0;
assign R3C34_GB30 = R3C33_GBO0;
assign R3C35_GB30 = R3C33_GBO0;
assign R3C32_GB30 = R3C33_GBO0;
assign R4C33_GB30 = R4C33_GBO0;
assign R4C34_GB30 = R4C33_GBO0;
assign R4C35_GB30 = R4C33_GBO0;
assign R4C32_GB30 = R4C33_GBO0;
assign R5C33_GB30 = R5C33_GBO0;
assign R5C34_GB30 = R5C33_GBO0;
assign R5C35_GB30 = R5C33_GBO0;
assign R5C32_GB30 = R5C33_GBO0;
assign R6C33_GB30 = R6C33_GBO0;
assign R6C34_GB30 = R6C33_GBO0;
assign R6C35_GB30 = R6C33_GBO0;
assign R6C32_GB30 = R6C33_GBO0;
assign R7C33_GB30 = R7C33_GBO0;
assign R7C34_GB30 = R7C33_GBO0;
assign R7C35_GB30 = R7C33_GBO0;
assign R7C32_GB30 = R7C33_GBO0;
assign R8C33_GB30 = R8C33_GBO0;
assign R8C34_GB30 = R8C33_GBO0;
assign R8C35_GB30 = R8C33_GBO0;
assign R8C32_GB30 = R8C33_GBO0;
assign R9C33_GB30 = R9C33_GBO0;
assign R9C34_GB30 = R9C33_GBO0;
assign R9C35_GB30 = R9C33_GBO0;
assign R9C32_GB30 = R9C33_GBO0;
assign R2C36_GB30 = R2C37_GBO0;
assign R2C37_GB30 = R2C37_GBO0;
assign R2C38_GB30 = R2C37_GBO0;
assign R2C39_GB30 = R2C37_GBO0;
assign R3C36_GB30 = R3C37_GBO0;
assign R3C37_GB30 = R3C37_GBO0;
assign R3C38_GB30 = R3C37_GBO0;
assign R3C39_GB30 = R3C37_GBO0;
assign R4C36_GB30 = R4C37_GBO0;
assign R4C37_GB30 = R4C37_GBO0;
assign R4C38_GB30 = R4C37_GBO0;
assign R4C39_GB30 = R4C37_GBO0;
assign R5C36_GB30 = R5C37_GBO0;
assign R5C37_GB30 = R5C37_GBO0;
assign R5C38_GB30 = R5C37_GBO0;
assign R5C39_GB30 = R5C37_GBO0;
assign R6C36_GB30 = R6C37_GBO0;
assign R6C37_GB30 = R6C37_GBO0;
assign R6C38_GB30 = R6C37_GBO0;
assign R6C39_GB30 = R6C37_GBO0;
assign R7C36_GB30 = R7C37_GBO0;
assign R7C37_GB30 = R7C37_GBO0;
assign R7C38_GB30 = R7C37_GBO0;
assign R7C39_GB30 = R7C37_GBO0;
assign R8C36_GB30 = R8C37_GBO0;
assign R8C37_GB30 = R8C37_GBO0;
assign R8C38_GB30 = R8C37_GBO0;
assign R8C39_GB30 = R8C37_GBO0;
assign R9C36_GB30 = R9C37_GBO0;
assign R9C37_GB30 = R9C37_GBO0;
assign R9C38_GB30 = R9C37_GBO0;
assign R9C39_GB30 = R9C37_GBO0;
assign R2C41_GB30 = R2C41_GBO0;
assign R2C42_GB30 = R2C41_GBO0;
assign R2C43_GB30 = R2C41_GBO0;
assign R2C40_GB30 = R2C41_GBO0;
assign R3C41_GB30 = R3C41_GBO0;
assign R3C42_GB30 = R3C41_GBO0;
assign R3C43_GB30 = R3C41_GBO0;
assign R3C40_GB30 = R3C41_GBO0;
assign R4C41_GB30 = R4C41_GBO0;
assign R4C42_GB30 = R4C41_GBO0;
assign R4C43_GB30 = R4C41_GBO0;
assign R4C40_GB30 = R4C41_GBO0;
assign R5C41_GB30 = R5C41_GBO0;
assign R5C42_GB30 = R5C41_GBO0;
assign R5C43_GB30 = R5C41_GBO0;
assign R5C40_GB30 = R5C41_GBO0;
assign R6C41_GB30 = R6C41_GBO0;
assign R6C42_GB30 = R6C41_GBO0;
assign R6C43_GB30 = R6C41_GBO0;
assign R6C40_GB30 = R6C41_GBO0;
assign R7C41_GB30 = R7C41_GBO0;
assign R7C42_GB30 = R7C41_GBO0;
assign R7C43_GB30 = R7C41_GBO0;
assign R7C40_GB30 = R7C41_GBO0;
assign R8C41_GB30 = R8C41_GBO0;
assign R8C42_GB30 = R8C41_GBO0;
assign R8C43_GB30 = R8C41_GBO0;
assign R8C40_GB30 = R8C41_GBO0;
assign R9C41_GB30 = R9C41_GBO0;
assign R9C42_GB30 = R9C41_GBO0;
assign R9C43_GB30 = R9C41_GBO0;
assign R9C40_GB30 = R9C41_GBO0;
assign R2C44_GB30 = R2C45_GBO0;
assign R2C45_GB30 = R2C45_GBO0;
assign R2C46_GB30 = R2C45_GBO0;
assign R3C44_GB30 = R3C45_GBO0;
assign R3C45_GB30 = R3C45_GBO0;
assign R3C46_GB30 = R3C45_GBO0;
assign R4C44_GB30 = R4C45_GBO0;
assign R4C45_GB30 = R4C45_GBO0;
assign R4C46_GB30 = R4C45_GBO0;
assign R5C44_GB30 = R5C45_GBO0;
assign R5C45_GB30 = R5C45_GBO0;
assign R5C46_GB30 = R5C45_GBO0;
assign R6C44_GB30 = R6C45_GBO0;
assign R6C45_GB30 = R6C45_GBO0;
assign R6C46_GB30 = R6C45_GBO0;
assign R7C44_GB30 = R7C45_GBO0;
assign R7C45_GB30 = R7C45_GBO0;
assign R7C46_GB30 = R7C45_GBO0;
assign R8C44_GB30 = R8C45_GBO0;
assign R8C45_GB30 = R8C45_GBO0;
assign R8C46_GB30 = R8C45_GBO0;
assign R9C44_GB30 = R9C45_GBO0;
assign R9C45_GB30 = R9C45_GBO0;
assign R9C46_GB30 = R9C45_GBO0;
assign R2C33_GB40 = R2C32_GBO1;
assign R2C34_GB40 = R2C32_GBO1;
assign R2C29_GB40 = R2C32_GBO1;
assign R2C30_GB40 = R2C32_GBO1;
assign R2C31_GB40 = R2C32_GBO1;
assign R2C32_GB40 = R2C32_GBO1;
assign R3C33_GB40 = R3C32_GBO1;
assign R3C34_GB40 = R3C32_GBO1;
assign R3C29_GB40 = R3C32_GBO1;
assign R3C30_GB40 = R3C32_GBO1;
assign R3C31_GB40 = R3C32_GBO1;
assign R3C32_GB40 = R3C32_GBO1;
assign R4C33_GB40 = R4C32_GBO1;
assign R4C34_GB40 = R4C32_GBO1;
assign R4C29_GB40 = R4C32_GBO1;
assign R4C30_GB40 = R4C32_GBO1;
assign R4C31_GB40 = R4C32_GBO1;
assign R4C32_GB40 = R4C32_GBO1;
assign R5C33_GB40 = R5C32_GBO1;
assign R5C34_GB40 = R5C32_GBO1;
assign R5C29_GB40 = R5C32_GBO1;
assign R5C30_GB40 = R5C32_GBO1;
assign R5C31_GB40 = R5C32_GBO1;
assign R5C32_GB40 = R5C32_GBO1;
assign R6C33_GB40 = R6C32_GBO1;
assign R6C34_GB40 = R6C32_GBO1;
assign R6C29_GB40 = R6C32_GBO1;
assign R6C30_GB40 = R6C32_GBO1;
assign R6C31_GB40 = R6C32_GBO1;
assign R6C32_GB40 = R6C32_GBO1;
assign R7C33_GB40 = R7C32_GBO1;
assign R7C34_GB40 = R7C32_GBO1;
assign R7C29_GB40 = R7C32_GBO1;
assign R7C30_GB40 = R7C32_GBO1;
assign R7C31_GB40 = R7C32_GBO1;
assign R7C32_GB40 = R7C32_GBO1;
assign R8C33_GB40 = R8C32_GBO1;
assign R8C34_GB40 = R8C32_GBO1;
assign R8C29_GB40 = R8C32_GBO1;
assign R8C30_GB40 = R8C32_GBO1;
assign R8C31_GB40 = R8C32_GBO1;
assign R8C32_GB40 = R8C32_GBO1;
assign R9C33_GB40 = R9C32_GBO1;
assign R9C34_GB40 = R9C32_GBO1;
assign R9C29_GB40 = R9C32_GBO1;
assign R9C30_GB40 = R9C32_GBO1;
assign R9C31_GB40 = R9C32_GBO1;
assign R9C32_GB40 = R9C32_GBO1;
assign R2C35_GB40 = R2C36_GBO1;
assign R2C36_GB40 = R2C36_GBO1;
assign R2C37_GB40 = R2C36_GBO1;
assign R2C38_GB40 = R2C36_GBO1;
assign R3C35_GB40 = R3C36_GBO1;
assign R3C36_GB40 = R3C36_GBO1;
assign R3C37_GB40 = R3C36_GBO1;
assign R3C38_GB40 = R3C36_GBO1;
assign R4C35_GB40 = R4C36_GBO1;
assign R4C36_GB40 = R4C36_GBO1;
assign R4C37_GB40 = R4C36_GBO1;
assign R4C38_GB40 = R4C36_GBO1;
assign R5C35_GB40 = R5C36_GBO1;
assign R5C36_GB40 = R5C36_GBO1;
assign R5C37_GB40 = R5C36_GBO1;
assign R5C38_GB40 = R5C36_GBO1;
assign R6C35_GB40 = R6C36_GBO1;
assign R6C36_GB40 = R6C36_GBO1;
assign R6C37_GB40 = R6C36_GBO1;
assign R6C38_GB40 = R6C36_GBO1;
assign R7C35_GB40 = R7C36_GBO1;
assign R7C36_GB40 = R7C36_GBO1;
assign R7C37_GB40 = R7C36_GBO1;
assign R7C38_GB40 = R7C36_GBO1;
assign R8C35_GB40 = R8C36_GBO1;
assign R8C36_GB40 = R8C36_GBO1;
assign R8C37_GB40 = R8C36_GBO1;
assign R8C38_GB40 = R8C36_GBO1;
assign R9C35_GB40 = R9C36_GBO1;
assign R9C36_GB40 = R9C36_GBO1;
assign R9C37_GB40 = R9C36_GBO1;
assign R9C38_GB40 = R9C36_GBO1;
assign R2C41_GB40 = R2C40_GBO1;
assign R2C42_GB40 = R2C40_GBO1;
assign R2C39_GB40 = R2C40_GBO1;
assign R2C40_GB40 = R2C40_GBO1;
assign R3C41_GB40 = R3C40_GBO1;
assign R3C42_GB40 = R3C40_GBO1;
assign R3C39_GB40 = R3C40_GBO1;
assign R3C40_GB40 = R3C40_GBO1;
assign R4C41_GB40 = R4C40_GBO1;
assign R4C42_GB40 = R4C40_GBO1;
assign R4C39_GB40 = R4C40_GBO1;
assign R4C40_GB40 = R4C40_GBO1;
assign R5C41_GB40 = R5C40_GBO1;
assign R5C42_GB40 = R5C40_GBO1;
assign R5C39_GB40 = R5C40_GBO1;
assign R5C40_GB40 = R5C40_GBO1;
assign R6C41_GB40 = R6C40_GBO1;
assign R6C42_GB40 = R6C40_GBO1;
assign R6C39_GB40 = R6C40_GBO1;
assign R6C40_GB40 = R6C40_GBO1;
assign R7C41_GB40 = R7C40_GBO1;
assign R7C42_GB40 = R7C40_GBO1;
assign R7C39_GB40 = R7C40_GBO1;
assign R7C40_GB40 = R7C40_GBO1;
assign R8C41_GB40 = R8C40_GBO1;
assign R8C42_GB40 = R8C40_GBO1;
assign R8C39_GB40 = R8C40_GBO1;
assign R8C40_GB40 = R8C40_GBO1;
assign R9C41_GB40 = R9C40_GBO1;
assign R9C42_GB40 = R9C40_GBO1;
assign R9C39_GB40 = R9C40_GBO1;
assign R9C40_GB40 = R9C40_GBO1;
assign R2C43_GB40 = R2C44_GBO1;
assign R2C44_GB40 = R2C44_GBO1;
assign R2C45_GB40 = R2C44_GBO1;
assign R2C46_GB40 = R2C44_GBO1;
assign R3C43_GB40 = R3C44_GBO1;
assign R3C44_GB40 = R3C44_GBO1;
assign R3C45_GB40 = R3C44_GBO1;
assign R3C46_GB40 = R3C44_GBO1;
assign R4C43_GB40 = R4C44_GBO1;
assign R4C44_GB40 = R4C44_GBO1;
assign R4C45_GB40 = R4C44_GBO1;
assign R4C46_GB40 = R4C44_GBO1;
assign R5C43_GB40 = R5C44_GBO1;
assign R5C44_GB40 = R5C44_GBO1;
assign R5C45_GB40 = R5C44_GBO1;
assign R5C46_GB40 = R5C44_GBO1;
assign R6C43_GB40 = R6C44_GBO1;
assign R6C44_GB40 = R6C44_GBO1;
assign R6C45_GB40 = R6C44_GBO1;
assign R6C46_GB40 = R6C44_GBO1;
assign R7C43_GB40 = R7C44_GBO1;
assign R7C44_GB40 = R7C44_GBO1;
assign R7C45_GB40 = R7C44_GBO1;
assign R7C46_GB40 = R7C44_GBO1;
assign R8C43_GB40 = R8C44_GBO1;
assign R8C44_GB40 = R8C44_GBO1;
assign R8C45_GB40 = R8C44_GBO1;
assign R8C46_GB40 = R8C44_GBO1;
assign R9C43_GB40 = R9C44_GBO1;
assign R9C44_GB40 = R9C44_GBO1;
assign R9C45_GB40 = R9C44_GBO1;
assign R9C46_GB40 = R9C44_GBO1;
assign R2C33_GB50 = R2C31_GBO1;
assign R2C29_GB50 = R2C31_GBO1;
assign R2C30_GB50 = R2C31_GBO1;
assign R2C31_GB50 = R2C31_GBO1;
assign R2C32_GB50 = R2C31_GBO1;
assign R3C33_GB50 = R3C31_GBO1;
assign R3C29_GB50 = R3C31_GBO1;
assign R3C30_GB50 = R3C31_GBO1;
assign R3C31_GB50 = R3C31_GBO1;
assign R3C32_GB50 = R3C31_GBO1;
assign R4C33_GB50 = R4C31_GBO1;
assign R4C29_GB50 = R4C31_GBO1;
assign R4C30_GB50 = R4C31_GBO1;
assign R4C31_GB50 = R4C31_GBO1;
assign R4C32_GB50 = R4C31_GBO1;
assign R5C33_GB50 = R5C31_GBO1;
assign R5C29_GB50 = R5C31_GBO1;
assign R5C30_GB50 = R5C31_GBO1;
assign R5C31_GB50 = R5C31_GBO1;
assign R5C32_GB50 = R5C31_GBO1;
assign R6C33_GB50 = R6C31_GBO1;
assign R6C29_GB50 = R6C31_GBO1;
assign R6C30_GB50 = R6C31_GBO1;
assign R6C31_GB50 = R6C31_GBO1;
assign R6C32_GB50 = R6C31_GBO1;
assign R7C33_GB50 = R7C31_GBO1;
assign R7C29_GB50 = R7C31_GBO1;
assign R7C30_GB50 = R7C31_GBO1;
assign R7C31_GB50 = R7C31_GBO1;
assign R7C32_GB50 = R7C31_GBO1;
assign R8C33_GB50 = R8C31_GBO1;
assign R8C29_GB50 = R8C31_GBO1;
assign R8C30_GB50 = R8C31_GBO1;
assign R8C31_GB50 = R8C31_GBO1;
assign R8C32_GB50 = R8C31_GBO1;
assign R9C33_GB50 = R9C31_GBO1;
assign R9C29_GB50 = R9C31_GBO1;
assign R9C30_GB50 = R9C31_GBO1;
assign R9C31_GB50 = R9C31_GBO1;
assign R9C32_GB50 = R9C31_GBO1;
assign R2C34_GB50 = R2C35_GBO1;
assign R2C35_GB50 = R2C35_GBO1;
assign R2C36_GB50 = R2C35_GBO1;
assign R2C37_GB50 = R2C35_GBO1;
assign R3C34_GB50 = R3C35_GBO1;
assign R3C35_GB50 = R3C35_GBO1;
assign R3C36_GB50 = R3C35_GBO1;
assign R3C37_GB50 = R3C35_GBO1;
assign R4C34_GB50 = R4C35_GBO1;
assign R4C35_GB50 = R4C35_GBO1;
assign R4C36_GB50 = R4C35_GBO1;
assign R4C37_GB50 = R4C35_GBO1;
assign R5C34_GB50 = R5C35_GBO1;
assign R5C35_GB50 = R5C35_GBO1;
assign R5C36_GB50 = R5C35_GBO1;
assign R5C37_GB50 = R5C35_GBO1;
assign R6C34_GB50 = R6C35_GBO1;
assign R6C35_GB50 = R6C35_GBO1;
assign R6C36_GB50 = R6C35_GBO1;
assign R6C37_GB50 = R6C35_GBO1;
assign R7C34_GB50 = R7C35_GBO1;
assign R7C35_GB50 = R7C35_GBO1;
assign R7C36_GB50 = R7C35_GBO1;
assign R7C37_GB50 = R7C35_GBO1;
assign R8C34_GB50 = R8C35_GBO1;
assign R8C35_GB50 = R8C35_GBO1;
assign R8C36_GB50 = R8C35_GBO1;
assign R8C37_GB50 = R8C35_GBO1;
assign R9C34_GB50 = R9C35_GBO1;
assign R9C35_GB50 = R9C35_GBO1;
assign R9C36_GB50 = R9C35_GBO1;
assign R9C37_GB50 = R9C35_GBO1;
assign R2C41_GB50 = R2C39_GBO1;
assign R2C38_GB50 = R2C39_GBO1;
assign R2C39_GB50 = R2C39_GBO1;
assign R2C40_GB50 = R2C39_GBO1;
assign R3C41_GB50 = R3C39_GBO1;
assign R3C38_GB50 = R3C39_GBO1;
assign R3C39_GB50 = R3C39_GBO1;
assign R3C40_GB50 = R3C39_GBO1;
assign R4C41_GB50 = R4C39_GBO1;
assign R4C38_GB50 = R4C39_GBO1;
assign R4C39_GB50 = R4C39_GBO1;
assign R4C40_GB50 = R4C39_GBO1;
assign R5C41_GB50 = R5C39_GBO1;
assign R5C38_GB50 = R5C39_GBO1;
assign R5C39_GB50 = R5C39_GBO1;
assign R5C40_GB50 = R5C39_GBO1;
assign R6C41_GB50 = R6C39_GBO1;
assign R6C38_GB50 = R6C39_GBO1;
assign R6C39_GB50 = R6C39_GBO1;
assign R6C40_GB50 = R6C39_GBO1;
assign R7C41_GB50 = R7C39_GBO1;
assign R7C38_GB50 = R7C39_GBO1;
assign R7C39_GB50 = R7C39_GBO1;
assign R7C40_GB50 = R7C39_GBO1;
assign R8C41_GB50 = R8C39_GBO1;
assign R8C38_GB50 = R8C39_GBO1;
assign R8C39_GB50 = R8C39_GBO1;
assign R8C40_GB50 = R8C39_GBO1;
assign R9C41_GB50 = R9C39_GBO1;
assign R9C38_GB50 = R9C39_GBO1;
assign R9C39_GB50 = R9C39_GBO1;
assign R9C40_GB50 = R9C39_GBO1;
assign R2C42_GB50 = R2C43_GBO1;
assign R2C43_GB50 = R2C43_GBO1;
assign R2C44_GB50 = R2C43_GBO1;
assign R2C45_GB50 = R2C43_GBO1;
assign R2C46_GB50 = R2C43_GBO1;
assign R3C42_GB50 = R3C43_GBO1;
assign R3C43_GB50 = R3C43_GBO1;
assign R3C44_GB50 = R3C43_GBO1;
assign R3C45_GB50 = R3C43_GBO1;
assign R3C46_GB50 = R3C43_GBO1;
assign R4C42_GB50 = R4C43_GBO1;
assign R4C43_GB50 = R4C43_GBO1;
assign R4C44_GB50 = R4C43_GBO1;
assign R4C45_GB50 = R4C43_GBO1;
assign R4C46_GB50 = R4C43_GBO1;
assign R5C42_GB50 = R5C43_GBO1;
assign R5C43_GB50 = R5C43_GBO1;
assign R5C44_GB50 = R5C43_GBO1;
assign R5C45_GB50 = R5C43_GBO1;
assign R5C46_GB50 = R5C43_GBO1;
assign R6C42_GB50 = R6C43_GBO1;
assign R6C43_GB50 = R6C43_GBO1;
assign R6C44_GB50 = R6C43_GBO1;
assign R6C45_GB50 = R6C43_GBO1;
assign R6C46_GB50 = R6C43_GBO1;
assign R7C42_GB50 = R7C43_GBO1;
assign R7C43_GB50 = R7C43_GBO1;
assign R7C44_GB50 = R7C43_GBO1;
assign R7C45_GB50 = R7C43_GBO1;
assign R7C46_GB50 = R7C43_GBO1;
assign R8C42_GB50 = R8C43_GBO1;
assign R8C43_GB50 = R8C43_GBO1;
assign R8C44_GB50 = R8C43_GBO1;
assign R8C45_GB50 = R8C43_GBO1;
assign R8C46_GB50 = R8C43_GBO1;
assign R9C42_GB50 = R9C43_GBO1;
assign R9C43_GB50 = R9C43_GBO1;
assign R9C44_GB50 = R9C43_GBO1;
assign R9C45_GB50 = R9C43_GBO1;
assign R9C46_GB50 = R9C43_GBO1;
assign R2C29_GB60 = R2C30_GBO1;
assign R2C30_GB60 = R2C30_GBO1;
assign R2C31_GB60 = R2C30_GBO1;
assign R2C32_GB60 = R2C30_GBO1;
assign R3C29_GB60 = R3C30_GBO1;
assign R3C30_GB60 = R3C30_GBO1;
assign R3C31_GB60 = R3C30_GBO1;
assign R3C32_GB60 = R3C30_GBO1;
assign R4C29_GB60 = R4C30_GBO1;
assign R4C30_GB60 = R4C30_GBO1;
assign R4C31_GB60 = R4C30_GBO1;
assign R4C32_GB60 = R4C30_GBO1;
assign R5C29_GB60 = R5C30_GBO1;
assign R5C30_GB60 = R5C30_GBO1;
assign R5C31_GB60 = R5C30_GBO1;
assign R5C32_GB60 = R5C30_GBO1;
assign R6C29_GB60 = R6C30_GBO1;
assign R6C30_GB60 = R6C30_GBO1;
assign R6C31_GB60 = R6C30_GBO1;
assign R6C32_GB60 = R6C30_GBO1;
assign R7C29_GB60 = R7C30_GBO1;
assign R7C30_GB60 = R7C30_GBO1;
assign R7C31_GB60 = R7C30_GBO1;
assign R7C32_GB60 = R7C30_GBO1;
assign R8C29_GB60 = R8C30_GBO1;
assign R8C30_GB60 = R8C30_GBO1;
assign R8C31_GB60 = R8C30_GBO1;
assign R8C32_GB60 = R8C30_GBO1;
assign R9C29_GB60 = R9C30_GBO1;
assign R9C30_GB60 = R9C30_GBO1;
assign R9C31_GB60 = R9C30_GBO1;
assign R9C32_GB60 = R9C30_GBO1;
assign R2C33_GB60 = R2C34_GBO1;
assign R2C34_GB60 = R2C34_GBO1;
assign R2C35_GB60 = R2C34_GBO1;
assign R2C36_GB60 = R2C34_GBO1;
assign R3C33_GB60 = R3C34_GBO1;
assign R3C34_GB60 = R3C34_GBO1;
assign R3C35_GB60 = R3C34_GBO1;
assign R3C36_GB60 = R3C34_GBO1;
assign R4C33_GB60 = R4C34_GBO1;
assign R4C34_GB60 = R4C34_GBO1;
assign R4C35_GB60 = R4C34_GBO1;
assign R4C36_GB60 = R4C34_GBO1;
assign R5C33_GB60 = R5C34_GBO1;
assign R5C34_GB60 = R5C34_GBO1;
assign R5C35_GB60 = R5C34_GBO1;
assign R5C36_GB60 = R5C34_GBO1;
assign R6C33_GB60 = R6C34_GBO1;
assign R6C34_GB60 = R6C34_GBO1;
assign R6C35_GB60 = R6C34_GBO1;
assign R6C36_GB60 = R6C34_GBO1;
assign R7C33_GB60 = R7C34_GBO1;
assign R7C34_GB60 = R7C34_GBO1;
assign R7C35_GB60 = R7C34_GBO1;
assign R7C36_GB60 = R7C34_GBO1;
assign R8C33_GB60 = R8C34_GBO1;
assign R8C34_GB60 = R8C34_GBO1;
assign R8C35_GB60 = R8C34_GBO1;
assign R8C36_GB60 = R8C34_GBO1;
assign R9C33_GB60 = R9C34_GBO1;
assign R9C34_GB60 = R9C34_GBO1;
assign R9C35_GB60 = R9C34_GBO1;
assign R9C36_GB60 = R9C34_GBO1;
assign R2C37_GB60 = R2C38_GBO1;
assign R2C38_GB60 = R2C38_GBO1;
assign R2C39_GB60 = R2C38_GBO1;
assign R2C40_GB60 = R2C38_GBO1;
assign R3C37_GB60 = R3C38_GBO1;
assign R3C38_GB60 = R3C38_GBO1;
assign R3C39_GB60 = R3C38_GBO1;
assign R3C40_GB60 = R3C38_GBO1;
assign R4C37_GB60 = R4C38_GBO1;
assign R4C38_GB60 = R4C38_GBO1;
assign R4C39_GB60 = R4C38_GBO1;
assign R4C40_GB60 = R4C38_GBO1;
assign R5C37_GB60 = R5C38_GBO1;
assign R5C38_GB60 = R5C38_GBO1;
assign R5C39_GB60 = R5C38_GBO1;
assign R5C40_GB60 = R5C38_GBO1;
assign R6C37_GB60 = R6C38_GBO1;
assign R6C38_GB60 = R6C38_GBO1;
assign R6C39_GB60 = R6C38_GBO1;
assign R6C40_GB60 = R6C38_GBO1;
assign R7C37_GB60 = R7C38_GBO1;
assign R7C38_GB60 = R7C38_GBO1;
assign R7C39_GB60 = R7C38_GBO1;
assign R7C40_GB60 = R7C38_GBO1;
assign R8C37_GB60 = R8C38_GBO1;
assign R8C38_GB60 = R8C38_GBO1;
assign R8C39_GB60 = R8C38_GBO1;
assign R8C40_GB60 = R8C38_GBO1;
assign R9C37_GB60 = R9C38_GBO1;
assign R9C38_GB60 = R9C38_GBO1;
assign R9C39_GB60 = R9C38_GBO1;
assign R9C40_GB60 = R9C38_GBO1;
assign R2C41_GB60 = R2C42_GBO1;
assign R2C42_GB60 = R2C42_GBO1;
assign R2C43_GB60 = R2C42_GBO1;
assign R2C44_GB60 = R2C42_GBO1;
assign R3C41_GB60 = R3C42_GBO1;
assign R3C42_GB60 = R3C42_GBO1;
assign R3C43_GB60 = R3C42_GBO1;
assign R3C44_GB60 = R3C42_GBO1;
assign R4C41_GB60 = R4C42_GBO1;
assign R4C42_GB60 = R4C42_GBO1;
assign R4C43_GB60 = R4C42_GBO1;
assign R4C44_GB60 = R4C42_GBO1;
assign R5C41_GB60 = R5C42_GBO1;
assign R5C42_GB60 = R5C42_GBO1;
assign R5C43_GB60 = R5C42_GBO1;
assign R5C44_GB60 = R5C42_GBO1;
assign R6C41_GB60 = R6C42_GBO1;
assign R6C42_GB60 = R6C42_GBO1;
assign R6C43_GB60 = R6C42_GBO1;
assign R6C44_GB60 = R6C42_GBO1;
assign R7C41_GB60 = R7C42_GBO1;
assign R7C42_GB60 = R7C42_GBO1;
assign R7C43_GB60 = R7C42_GBO1;
assign R7C44_GB60 = R7C42_GBO1;
assign R8C41_GB60 = R8C42_GBO1;
assign R8C42_GB60 = R8C42_GBO1;
assign R8C43_GB60 = R8C42_GBO1;
assign R8C44_GB60 = R8C42_GBO1;
assign R9C41_GB60 = R9C42_GBO1;
assign R9C42_GB60 = R9C42_GBO1;
assign R9C43_GB60 = R9C42_GBO1;
assign R9C44_GB60 = R9C42_GBO1;
assign R2C45_GB60 = R2C46_GBO1;
assign R2C46_GB60 = R2C46_GBO1;
assign R3C45_GB60 = R3C46_GBO1;
assign R3C46_GB60 = R3C46_GBO1;
assign R4C45_GB60 = R4C46_GBO1;
assign R4C46_GB60 = R4C46_GBO1;
assign R5C45_GB60 = R5C46_GBO1;
assign R5C46_GB60 = R5C46_GBO1;
assign R6C45_GB60 = R6C46_GBO1;
assign R6C46_GB60 = R6C46_GBO1;
assign R7C45_GB60 = R7C46_GBO1;
assign R7C46_GB60 = R7C46_GBO1;
assign R8C45_GB60 = R8C46_GBO1;
assign R8C46_GB60 = R8C46_GBO1;
assign R9C45_GB60 = R9C46_GBO1;
assign R9C46_GB60 = R9C46_GBO1;
assign R2C29_GB70 = R2C29_GBO1;
assign R2C30_GB70 = R2C29_GBO1;
assign R2C31_GB70 = R2C29_GBO1;
assign R3C29_GB70 = R3C29_GBO1;
assign R3C30_GB70 = R3C29_GBO1;
assign R3C31_GB70 = R3C29_GBO1;
assign R4C29_GB70 = R4C29_GBO1;
assign R4C30_GB70 = R4C29_GBO1;
assign R4C31_GB70 = R4C29_GBO1;
assign R5C29_GB70 = R5C29_GBO1;
assign R5C30_GB70 = R5C29_GBO1;
assign R5C31_GB70 = R5C29_GBO1;
assign R6C29_GB70 = R6C29_GBO1;
assign R6C30_GB70 = R6C29_GBO1;
assign R6C31_GB70 = R6C29_GBO1;
assign R7C29_GB70 = R7C29_GBO1;
assign R7C30_GB70 = R7C29_GBO1;
assign R7C31_GB70 = R7C29_GBO1;
assign R8C29_GB70 = R8C29_GBO1;
assign R8C30_GB70 = R8C29_GBO1;
assign R8C31_GB70 = R8C29_GBO1;
assign R9C29_GB70 = R9C29_GBO1;
assign R9C30_GB70 = R9C29_GBO1;
assign R9C31_GB70 = R9C29_GBO1;
assign R2C33_GB70 = R2C33_GBO1;
assign R2C34_GB70 = R2C33_GBO1;
assign R2C35_GB70 = R2C33_GBO1;
assign R2C32_GB70 = R2C33_GBO1;
assign R3C33_GB70 = R3C33_GBO1;
assign R3C34_GB70 = R3C33_GBO1;
assign R3C35_GB70 = R3C33_GBO1;
assign R3C32_GB70 = R3C33_GBO1;
assign R4C33_GB70 = R4C33_GBO1;
assign R4C34_GB70 = R4C33_GBO1;
assign R4C35_GB70 = R4C33_GBO1;
assign R4C32_GB70 = R4C33_GBO1;
assign R5C33_GB70 = R5C33_GBO1;
assign R5C34_GB70 = R5C33_GBO1;
assign R5C35_GB70 = R5C33_GBO1;
assign R5C32_GB70 = R5C33_GBO1;
assign R6C33_GB70 = R6C33_GBO1;
assign R6C34_GB70 = R6C33_GBO1;
assign R6C35_GB70 = R6C33_GBO1;
assign R6C32_GB70 = R6C33_GBO1;
assign R7C33_GB70 = R7C33_GBO1;
assign R7C34_GB70 = R7C33_GBO1;
assign R7C35_GB70 = R7C33_GBO1;
assign R7C32_GB70 = R7C33_GBO1;
assign R8C33_GB70 = R8C33_GBO1;
assign R8C34_GB70 = R8C33_GBO1;
assign R8C35_GB70 = R8C33_GBO1;
assign R8C32_GB70 = R8C33_GBO1;
assign R9C33_GB70 = R9C33_GBO1;
assign R9C34_GB70 = R9C33_GBO1;
assign R9C35_GB70 = R9C33_GBO1;
assign R9C32_GB70 = R9C33_GBO1;
assign R2C36_GB70 = R2C37_GBO1;
assign R2C37_GB70 = R2C37_GBO1;
assign R2C38_GB70 = R2C37_GBO1;
assign R2C39_GB70 = R2C37_GBO1;
assign R3C36_GB70 = R3C37_GBO1;
assign R3C37_GB70 = R3C37_GBO1;
assign R3C38_GB70 = R3C37_GBO1;
assign R3C39_GB70 = R3C37_GBO1;
assign R4C36_GB70 = R4C37_GBO1;
assign R4C37_GB70 = R4C37_GBO1;
assign R4C38_GB70 = R4C37_GBO1;
assign R4C39_GB70 = R4C37_GBO1;
assign R5C36_GB70 = R5C37_GBO1;
assign R5C37_GB70 = R5C37_GBO1;
assign R5C38_GB70 = R5C37_GBO1;
assign R5C39_GB70 = R5C37_GBO1;
assign R6C36_GB70 = R6C37_GBO1;
assign R6C37_GB70 = R6C37_GBO1;
assign R6C38_GB70 = R6C37_GBO1;
assign R6C39_GB70 = R6C37_GBO1;
assign R7C36_GB70 = R7C37_GBO1;
assign R7C37_GB70 = R7C37_GBO1;
assign R7C38_GB70 = R7C37_GBO1;
assign R7C39_GB70 = R7C37_GBO1;
assign R8C36_GB70 = R8C37_GBO1;
assign R8C37_GB70 = R8C37_GBO1;
assign R8C38_GB70 = R8C37_GBO1;
assign R8C39_GB70 = R8C37_GBO1;
assign R9C36_GB70 = R9C37_GBO1;
assign R9C37_GB70 = R9C37_GBO1;
assign R9C38_GB70 = R9C37_GBO1;
assign R9C39_GB70 = R9C37_GBO1;
assign R2C41_GB70 = R2C41_GBO1;
assign R2C42_GB70 = R2C41_GBO1;
assign R2C43_GB70 = R2C41_GBO1;
assign R2C40_GB70 = R2C41_GBO1;
assign R3C41_GB70 = R3C41_GBO1;
assign R3C42_GB70 = R3C41_GBO1;
assign R3C43_GB70 = R3C41_GBO1;
assign R3C40_GB70 = R3C41_GBO1;
assign R4C41_GB70 = R4C41_GBO1;
assign R4C42_GB70 = R4C41_GBO1;
assign R4C43_GB70 = R4C41_GBO1;
assign R4C40_GB70 = R4C41_GBO1;
assign R5C41_GB70 = R5C41_GBO1;
assign R5C42_GB70 = R5C41_GBO1;
assign R5C43_GB70 = R5C41_GBO1;
assign R5C40_GB70 = R5C41_GBO1;
assign R6C41_GB70 = R6C41_GBO1;
assign R6C42_GB70 = R6C41_GBO1;
assign R6C43_GB70 = R6C41_GBO1;
assign R6C40_GB70 = R6C41_GBO1;
assign R7C41_GB70 = R7C41_GBO1;
assign R7C42_GB70 = R7C41_GBO1;
assign R7C43_GB70 = R7C41_GBO1;
assign R7C40_GB70 = R7C41_GBO1;
assign R8C41_GB70 = R8C41_GBO1;
assign R8C42_GB70 = R8C41_GBO1;
assign R8C43_GB70 = R8C41_GBO1;
assign R8C40_GB70 = R8C41_GBO1;
assign R9C41_GB70 = R9C41_GBO1;
assign R9C42_GB70 = R9C41_GBO1;
assign R9C43_GB70 = R9C41_GBO1;
assign R9C40_GB70 = R9C41_GBO1;
assign R2C44_GB70 = R2C45_GBO1;
assign R2C45_GB70 = R2C45_GBO1;
assign R2C46_GB70 = R2C45_GBO1;
assign R3C44_GB70 = R3C45_GBO1;
assign R3C45_GB70 = R3C45_GBO1;
assign R3C46_GB70 = R3C45_GBO1;
assign R4C44_GB70 = R4C45_GBO1;
assign R4C45_GB70 = R4C45_GBO1;
assign R4C46_GB70 = R4C45_GBO1;
assign R5C44_GB70 = R5C45_GBO1;
assign R5C45_GB70 = R5C45_GBO1;
assign R5C46_GB70 = R5C45_GBO1;
assign R6C44_GB70 = R6C45_GBO1;
assign R6C45_GB70 = R6C45_GBO1;
assign R6C46_GB70 = R6C45_GBO1;
assign R7C44_GB70 = R7C45_GBO1;
assign R7C45_GB70 = R7C45_GBO1;
assign R7C46_GB70 = R7C45_GBO1;
assign R8C44_GB70 = R8C45_GBO1;
assign R8C45_GB70 = R8C45_GBO1;
assign R8C46_GB70 = R8C45_GBO1;
assign R9C44_GB70 = R9C45_GBO1;
assign R9C45_GB70 = R9C45_GBO1;
assign R9C46_GB70 = R9C45_GBO1;
assign R11C33_GB00 = R11C32_GBO0;
assign R11C34_GB00 = R11C32_GBO0;
assign R11C29_GB00 = R11C32_GBO0;
assign R11C30_GB00 = R11C32_GBO0;
assign R11C31_GB00 = R11C32_GBO0;
assign R11C32_GB00 = R11C32_GBO0;
assign R12C33_GB00 = R12C32_GBO0;
assign R12C34_GB00 = R12C32_GBO0;
assign R12C29_GB00 = R12C32_GBO0;
assign R12C30_GB00 = R12C32_GBO0;
assign R12C31_GB00 = R12C32_GBO0;
assign R12C32_GB00 = R12C32_GBO0;
assign R13C33_GB00 = R13C32_GBO0;
assign R13C34_GB00 = R13C32_GBO0;
assign R13C29_GB00 = R13C32_GBO0;
assign R13C30_GB00 = R13C32_GBO0;
assign R13C31_GB00 = R13C32_GBO0;
assign R13C32_GB00 = R13C32_GBO0;
assign R14C33_GB00 = R14C32_GBO0;
assign R14C34_GB00 = R14C32_GBO0;
assign R14C29_GB00 = R14C32_GBO0;
assign R14C30_GB00 = R14C32_GBO0;
assign R14C31_GB00 = R14C32_GBO0;
assign R14C32_GB00 = R14C32_GBO0;
assign R15C33_GB00 = R15C32_GBO0;
assign R15C34_GB00 = R15C32_GBO0;
assign R15C29_GB00 = R15C32_GBO0;
assign R15C30_GB00 = R15C32_GBO0;
assign R15C31_GB00 = R15C32_GBO0;
assign R15C32_GB00 = R15C32_GBO0;
assign R16C33_GB00 = R16C32_GBO0;
assign R16C34_GB00 = R16C32_GBO0;
assign R16C29_GB00 = R16C32_GBO0;
assign R16C30_GB00 = R16C32_GBO0;
assign R16C31_GB00 = R16C32_GBO0;
assign R16C32_GB00 = R16C32_GBO0;
assign R17C33_GB00 = R17C32_GBO0;
assign R17C34_GB00 = R17C32_GBO0;
assign R17C29_GB00 = R17C32_GBO0;
assign R17C30_GB00 = R17C32_GBO0;
assign R17C31_GB00 = R17C32_GBO0;
assign R17C32_GB00 = R17C32_GBO0;
assign R18C33_GB00 = R18C32_GBO0;
assign R18C34_GB00 = R18C32_GBO0;
assign R18C29_GB00 = R18C32_GBO0;
assign R18C30_GB00 = R18C32_GBO0;
assign R18C31_GB00 = R18C32_GBO0;
assign R18C32_GB00 = R18C32_GBO0;
assign R20C33_GB00 = R20C32_GBO0;
assign R20C34_GB00 = R20C32_GBO0;
assign R20C29_GB00 = R20C32_GBO0;
assign R20C30_GB00 = R20C32_GBO0;
assign R20C31_GB00 = R20C32_GBO0;
assign R20C32_GB00 = R20C32_GBO0;
assign R21C33_GB00 = R21C32_GBO0;
assign R21C34_GB00 = R21C32_GBO0;
assign R21C29_GB00 = R21C32_GBO0;
assign R21C30_GB00 = R21C32_GBO0;
assign R21C31_GB00 = R21C32_GBO0;
assign R21C32_GB00 = R21C32_GBO0;
assign R22C33_GB00 = R22C32_GBO0;
assign R22C34_GB00 = R22C32_GBO0;
assign R22C29_GB00 = R22C32_GBO0;
assign R22C30_GB00 = R22C32_GBO0;
assign R22C31_GB00 = R22C32_GBO0;
assign R22C32_GB00 = R22C32_GBO0;
assign R23C33_GB00 = R23C32_GBO0;
assign R23C34_GB00 = R23C32_GBO0;
assign R23C29_GB00 = R23C32_GBO0;
assign R23C30_GB00 = R23C32_GBO0;
assign R23C31_GB00 = R23C32_GBO0;
assign R23C32_GB00 = R23C32_GBO0;
assign R24C33_GB00 = R24C32_GBO0;
assign R24C34_GB00 = R24C32_GBO0;
assign R24C29_GB00 = R24C32_GBO0;
assign R24C30_GB00 = R24C32_GBO0;
assign R24C31_GB00 = R24C32_GBO0;
assign R24C32_GB00 = R24C32_GBO0;
assign R25C33_GB00 = R25C32_GBO0;
assign R25C34_GB00 = R25C32_GBO0;
assign R25C29_GB00 = R25C32_GBO0;
assign R25C30_GB00 = R25C32_GBO0;
assign R25C31_GB00 = R25C32_GBO0;
assign R25C32_GB00 = R25C32_GBO0;
assign R26C33_GB00 = R26C32_GBO0;
assign R26C34_GB00 = R26C32_GBO0;
assign R26C29_GB00 = R26C32_GBO0;
assign R26C30_GB00 = R26C32_GBO0;
assign R26C31_GB00 = R26C32_GBO0;
assign R26C32_GB00 = R26C32_GBO0;
assign R27C33_GB00 = R27C32_GBO0;
assign R27C34_GB00 = R27C32_GBO0;
assign R27C29_GB00 = R27C32_GBO0;
assign R27C30_GB00 = R27C32_GBO0;
assign R27C31_GB00 = R27C32_GBO0;
assign R27C32_GB00 = R27C32_GBO0;
assign R11C35_GB00 = R11C36_GBO0;
assign R11C36_GB00 = R11C36_GBO0;
assign R11C37_GB00 = R11C36_GBO0;
assign R11C38_GB00 = R11C36_GBO0;
assign R12C35_GB00 = R12C36_GBO0;
assign R12C36_GB00 = R12C36_GBO0;
assign R12C37_GB00 = R12C36_GBO0;
assign R12C38_GB00 = R12C36_GBO0;
assign R13C35_GB00 = R13C36_GBO0;
assign R13C36_GB00 = R13C36_GBO0;
assign R13C37_GB00 = R13C36_GBO0;
assign R13C38_GB00 = R13C36_GBO0;
assign R14C35_GB00 = R14C36_GBO0;
assign R14C36_GB00 = R14C36_GBO0;
assign R14C37_GB00 = R14C36_GBO0;
assign R14C38_GB00 = R14C36_GBO0;
assign R15C35_GB00 = R15C36_GBO0;
assign R15C36_GB00 = R15C36_GBO0;
assign R15C37_GB00 = R15C36_GBO0;
assign R15C38_GB00 = R15C36_GBO0;
assign R16C35_GB00 = R16C36_GBO0;
assign R16C36_GB00 = R16C36_GBO0;
assign R16C37_GB00 = R16C36_GBO0;
assign R16C38_GB00 = R16C36_GBO0;
assign R17C35_GB00 = R17C36_GBO0;
assign R17C36_GB00 = R17C36_GBO0;
assign R17C37_GB00 = R17C36_GBO0;
assign R17C38_GB00 = R17C36_GBO0;
assign R18C35_GB00 = R18C36_GBO0;
assign R18C36_GB00 = R18C36_GBO0;
assign R18C37_GB00 = R18C36_GBO0;
assign R18C38_GB00 = R18C36_GBO0;
assign R20C35_GB00 = R20C36_GBO0;
assign R20C36_GB00 = R20C36_GBO0;
assign R20C37_GB00 = R20C36_GBO0;
assign R20C38_GB00 = R20C36_GBO0;
assign R21C35_GB00 = R21C36_GBO0;
assign R21C36_GB00 = R21C36_GBO0;
assign R21C37_GB00 = R21C36_GBO0;
assign R21C38_GB00 = R21C36_GBO0;
assign R22C35_GB00 = R22C36_GBO0;
assign R22C36_GB00 = R22C36_GBO0;
assign R22C37_GB00 = R22C36_GBO0;
assign R22C38_GB00 = R22C36_GBO0;
assign R23C35_GB00 = R23C36_GBO0;
assign R23C36_GB00 = R23C36_GBO0;
assign R23C37_GB00 = R23C36_GBO0;
assign R23C38_GB00 = R23C36_GBO0;
assign R24C35_GB00 = R24C36_GBO0;
assign R24C36_GB00 = R24C36_GBO0;
assign R24C37_GB00 = R24C36_GBO0;
assign R24C38_GB00 = R24C36_GBO0;
assign R25C35_GB00 = R25C36_GBO0;
assign R25C36_GB00 = R25C36_GBO0;
assign R25C37_GB00 = R25C36_GBO0;
assign R25C38_GB00 = R25C36_GBO0;
assign R26C35_GB00 = R26C36_GBO0;
assign R26C36_GB00 = R26C36_GBO0;
assign R26C37_GB00 = R26C36_GBO0;
assign R26C38_GB00 = R26C36_GBO0;
assign R27C35_GB00 = R27C36_GBO0;
assign R27C36_GB00 = R27C36_GBO0;
assign R27C37_GB00 = R27C36_GBO0;
assign R27C38_GB00 = R27C36_GBO0;
assign R11C41_GB00 = R11C40_GBO0;
assign R11C42_GB00 = R11C40_GBO0;
assign R11C39_GB00 = R11C40_GBO0;
assign R11C40_GB00 = R11C40_GBO0;
assign R12C41_GB00 = R12C40_GBO0;
assign R12C42_GB00 = R12C40_GBO0;
assign R12C39_GB00 = R12C40_GBO0;
assign R12C40_GB00 = R12C40_GBO0;
assign R13C41_GB00 = R13C40_GBO0;
assign R13C42_GB00 = R13C40_GBO0;
assign R13C39_GB00 = R13C40_GBO0;
assign R13C40_GB00 = R13C40_GBO0;
assign R14C41_GB00 = R14C40_GBO0;
assign R14C42_GB00 = R14C40_GBO0;
assign R14C39_GB00 = R14C40_GBO0;
assign R14C40_GB00 = R14C40_GBO0;
assign R15C41_GB00 = R15C40_GBO0;
assign R15C42_GB00 = R15C40_GBO0;
assign R15C39_GB00 = R15C40_GBO0;
assign R15C40_GB00 = R15C40_GBO0;
assign R16C41_GB00 = R16C40_GBO0;
assign R16C42_GB00 = R16C40_GBO0;
assign R16C39_GB00 = R16C40_GBO0;
assign R16C40_GB00 = R16C40_GBO0;
assign R17C41_GB00 = R17C40_GBO0;
assign R17C42_GB00 = R17C40_GBO0;
assign R17C39_GB00 = R17C40_GBO0;
assign R17C40_GB00 = R17C40_GBO0;
assign R18C41_GB00 = R18C40_GBO0;
assign R18C42_GB00 = R18C40_GBO0;
assign R18C39_GB00 = R18C40_GBO0;
assign R18C40_GB00 = R18C40_GBO0;
assign R20C41_GB00 = R20C40_GBO0;
assign R20C42_GB00 = R20C40_GBO0;
assign R20C39_GB00 = R20C40_GBO0;
assign R20C40_GB00 = R20C40_GBO0;
assign R21C41_GB00 = R21C40_GBO0;
assign R21C42_GB00 = R21C40_GBO0;
assign R21C39_GB00 = R21C40_GBO0;
assign R21C40_GB00 = R21C40_GBO0;
assign R22C41_GB00 = R22C40_GBO0;
assign R22C42_GB00 = R22C40_GBO0;
assign R22C39_GB00 = R22C40_GBO0;
assign R22C40_GB00 = R22C40_GBO0;
assign R23C41_GB00 = R23C40_GBO0;
assign R23C42_GB00 = R23C40_GBO0;
assign R23C39_GB00 = R23C40_GBO0;
assign R23C40_GB00 = R23C40_GBO0;
assign R24C41_GB00 = R24C40_GBO0;
assign R24C42_GB00 = R24C40_GBO0;
assign R24C39_GB00 = R24C40_GBO0;
assign R24C40_GB00 = R24C40_GBO0;
assign R25C41_GB00 = R25C40_GBO0;
assign R25C42_GB00 = R25C40_GBO0;
assign R25C39_GB00 = R25C40_GBO0;
assign R25C40_GB00 = R25C40_GBO0;
assign R26C41_GB00 = R26C40_GBO0;
assign R26C42_GB00 = R26C40_GBO0;
assign R26C39_GB00 = R26C40_GBO0;
assign R26C40_GB00 = R26C40_GBO0;
assign R27C41_GB00 = R27C40_GBO0;
assign R27C42_GB00 = R27C40_GBO0;
assign R27C39_GB00 = R27C40_GBO0;
assign R27C40_GB00 = R27C40_GBO0;
assign R11C43_GB00 = R11C44_GBO0;
assign R11C44_GB00 = R11C44_GBO0;
assign R11C45_GB00 = R11C44_GBO0;
assign R11C46_GB00 = R11C44_GBO0;
assign R12C43_GB00 = R12C44_GBO0;
assign R12C44_GB00 = R12C44_GBO0;
assign R12C45_GB00 = R12C44_GBO0;
assign R12C46_GB00 = R12C44_GBO0;
assign R13C43_GB00 = R13C44_GBO0;
assign R13C44_GB00 = R13C44_GBO0;
assign R13C45_GB00 = R13C44_GBO0;
assign R13C46_GB00 = R13C44_GBO0;
assign R14C43_GB00 = R14C44_GBO0;
assign R14C44_GB00 = R14C44_GBO0;
assign R14C45_GB00 = R14C44_GBO0;
assign R14C46_GB00 = R14C44_GBO0;
assign R15C43_GB00 = R15C44_GBO0;
assign R15C44_GB00 = R15C44_GBO0;
assign R15C45_GB00 = R15C44_GBO0;
assign R15C46_GB00 = R15C44_GBO0;
assign R16C43_GB00 = R16C44_GBO0;
assign R16C44_GB00 = R16C44_GBO0;
assign R16C45_GB00 = R16C44_GBO0;
assign R16C46_GB00 = R16C44_GBO0;
assign R17C43_GB00 = R17C44_GBO0;
assign R17C44_GB00 = R17C44_GBO0;
assign R17C45_GB00 = R17C44_GBO0;
assign R17C46_GB00 = R17C44_GBO0;
assign R18C43_GB00 = R18C44_GBO0;
assign R18C44_GB00 = R18C44_GBO0;
assign R18C45_GB00 = R18C44_GBO0;
assign R18C46_GB00 = R18C44_GBO0;
assign R20C43_GB00 = R20C44_GBO0;
assign R20C44_GB00 = R20C44_GBO0;
assign R20C45_GB00 = R20C44_GBO0;
assign R20C46_GB00 = R20C44_GBO0;
assign R21C43_GB00 = R21C44_GBO0;
assign R21C44_GB00 = R21C44_GBO0;
assign R21C45_GB00 = R21C44_GBO0;
assign R21C46_GB00 = R21C44_GBO0;
assign R22C43_GB00 = R22C44_GBO0;
assign R22C44_GB00 = R22C44_GBO0;
assign R22C45_GB00 = R22C44_GBO0;
assign R22C46_GB00 = R22C44_GBO0;
assign R23C43_GB00 = R23C44_GBO0;
assign R23C44_GB00 = R23C44_GBO0;
assign R23C45_GB00 = R23C44_GBO0;
assign R23C46_GB00 = R23C44_GBO0;
assign R24C43_GB00 = R24C44_GBO0;
assign R24C44_GB00 = R24C44_GBO0;
assign R24C45_GB00 = R24C44_GBO0;
assign R24C46_GB00 = R24C44_GBO0;
assign R25C43_GB00 = R25C44_GBO0;
assign R25C44_GB00 = R25C44_GBO0;
assign R25C45_GB00 = R25C44_GBO0;
assign R25C46_GB00 = R25C44_GBO0;
assign R26C43_GB00 = R26C44_GBO0;
assign R26C44_GB00 = R26C44_GBO0;
assign R26C45_GB00 = R26C44_GBO0;
assign R26C46_GB00 = R26C44_GBO0;
assign R27C43_GB00 = R27C44_GBO0;
assign R27C44_GB00 = R27C44_GBO0;
assign R27C45_GB00 = R27C44_GBO0;
assign R27C46_GB00 = R27C44_GBO0;
assign R11C33_GB10 = R11C31_GBO0;
assign R11C29_GB10 = R11C31_GBO0;
assign R11C30_GB10 = R11C31_GBO0;
assign R11C31_GB10 = R11C31_GBO0;
assign R11C32_GB10 = R11C31_GBO0;
assign R12C33_GB10 = R12C31_GBO0;
assign R12C29_GB10 = R12C31_GBO0;
assign R12C30_GB10 = R12C31_GBO0;
assign R12C31_GB10 = R12C31_GBO0;
assign R12C32_GB10 = R12C31_GBO0;
assign R13C33_GB10 = R13C31_GBO0;
assign R13C29_GB10 = R13C31_GBO0;
assign R13C30_GB10 = R13C31_GBO0;
assign R13C31_GB10 = R13C31_GBO0;
assign R13C32_GB10 = R13C31_GBO0;
assign R14C33_GB10 = R14C31_GBO0;
assign R14C29_GB10 = R14C31_GBO0;
assign R14C30_GB10 = R14C31_GBO0;
assign R14C31_GB10 = R14C31_GBO0;
assign R14C32_GB10 = R14C31_GBO0;
assign R15C33_GB10 = R15C31_GBO0;
assign R15C29_GB10 = R15C31_GBO0;
assign R15C30_GB10 = R15C31_GBO0;
assign R15C31_GB10 = R15C31_GBO0;
assign R15C32_GB10 = R15C31_GBO0;
assign R16C33_GB10 = R16C31_GBO0;
assign R16C29_GB10 = R16C31_GBO0;
assign R16C30_GB10 = R16C31_GBO0;
assign R16C31_GB10 = R16C31_GBO0;
assign R16C32_GB10 = R16C31_GBO0;
assign R17C33_GB10 = R17C31_GBO0;
assign R17C29_GB10 = R17C31_GBO0;
assign R17C30_GB10 = R17C31_GBO0;
assign R17C31_GB10 = R17C31_GBO0;
assign R17C32_GB10 = R17C31_GBO0;
assign R18C33_GB10 = R18C31_GBO0;
assign R18C29_GB10 = R18C31_GBO0;
assign R18C30_GB10 = R18C31_GBO0;
assign R18C31_GB10 = R18C31_GBO0;
assign R18C32_GB10 = R18C31_GBO0;
assign R20C33_GB10 = R20C31_GBO0;
assign R20C29_GB10 = R20C31_GBO0;
assign R20C30_GB10 = R20C31_GBO0;
assign R20C31_GB10 = R20C31_GBO0;
assign R20C32_GB10 = R20C31_GBO0;
assign R21C33_GB10 = R21C31_GBO0;
assign R21C29_GB10 = R21C31_GBO0;
assign R21C30_GB10 = R21C31_GBO0;
assign R21C31_GB10 = R21C31_GBO0;
assign R21C32_GB10 = R21C31_GBO0;
assign R22C33_GB10 = R22C31_GBO0;
assign R22C29_GB10 = R22C31_GBO0;
assign R22C30_GB10 = R22C31_GBO0;
assign R22C31_GB10 = R22C31_GBO0;
assign R22C32_GB10 = R22C31_GBO0;
assign R23C33_GB10 = R23C31_GBO0;
assign R23C29_GB10 = R23C31_GBO0;
assign R23C30_GB10 = R23C31_GBO0;
assign R23C31_GB10 = R23C31_GBO0;
assign R23C32_GB10 = R23C31_GBO0;
assign R24C33_GB10 = R24C31_GBO0;
assign R24C29_GB10 = R24C31_GBO0;
assign R24C30_GB10 = R24C31_GBO0;
assign R24C31_GB10 = R24C31_GBO0;
assign R24C32_GB10 = R24C31_GBO0;
assign R25C33_GB10 = R25C31_GBO0;
assign R25C29_GB10 = R25C31_GBO0;
assign R25C30_GB10 = R25C31_GBO0;
assign R25C31_GB10 = R25C31_GBO0;
assign R25C32_GB10 = R25C31_GBO0;
assign R26C33_GB10 = R26C31_GBO0;
assign R26C29_GB10 = R26C31_GBO0;
assign R26C30_GB10 = R26C31_GBO0;
assign R26C31_GB10 = R26C31_GBO0;
assign R26C32_GB10 = R26C31_GBO0;
assign R27C33_GB10 = R27C31_GBO0;
assign R27C29_GB10 = R27C31_GBO0;
assign R27C30_GB10 = R27C31_GBO0;
assign R27C31_GB10 = R27C31_GBO0;
assign R27C32_GB10 = R27C31_GBO0;
assign R11C34_GB10 = R11C35_GBO0;
assign R11C35_GB10 = R11C35_GBO0;
assign R11C36_GB10 = R11C35_GBO0;
assign R11C37_GB10 = R11C35_GBO0;
assign R12C34_GB10 = R12C35_GBO0;
assign R12C35_GB10 = R12C35_GBO0;
assign R12C36_GB10 = R12C35_GBO0;
assign R12C37_GB10 = R12C35_GBO0;
assign R13C34_GB10 = R13C35_GBO0;
assign R13C35_GB10 = R13C35_GBO0;
assign R13C36_GB10 = R13C35_GBO0;
assign R13C37_GB10 = R13C35_GBO0;
assign R14C34_GB10 = R14C35_GBO0;
assign R14C35_GB10 = R14C35_GBO0;
assign R14C36_GB10 = R14C35_GBO0;
assign R14C37_GB10 = R14C35_GBO0;
assign R15C34_GB10 = R15C35_GBO0;
assign R15C35_GB10 = R15C35_GBO0;
assign R15C36_GB10 = R15C35_GBO0;
assign R15C37_GB10 = R15C35_GBO0;
assign R16C34_GB10 = R16C35_GBO0;
assign R16C35_GB10 = R16C35_GBO0;
assign R16C36_GB10 = R16C35_GBO0;
assign R16C37_GB10 = R16C35_GBO0;
assign R17C34_GB10 = R17C35_GBO0;
assign R17C35_GB10 = R17C35_GBO0;
assign R17C36_GB10 = R17C35_GBO0;
assign R17C37_GB10 = R17C35_GBO0;
assign R18C34_GB10 = R18C35_GBO0;
assign R18C35_GB10 = R18C35_GBO0;
assign R18C36_GB10 = R18C35_GBO0;
assign R18C37_GB10 = R18C35_GBO0;
assign R20C34_GB10 = R20C35_GBO0;
assign R20C35_GB10 = R20C35_GBO0;
assign R20C36_GB10 = R20C35_GBO0;
assign R20C37_GB10 = R20C35_GBO0;
assign R21C34_GB10 = R21C35_GBO0;
assign R21C35_GB10 = R21C35_GBO0;
assign R21C36_GB10 = R21C35_GBO0;
assign R21C37_GB10 = R21C35_GBO0;
assign R22C34_GB10 = R22C35_GBO0;
assign R22C35_GB10 = R22C35_GBO0;
assign R22C36_GB10 = R22C35_GBO0;
assign R22C37_GB10 = R22C35_GBO0;
assign R23C34_GB10 = R23C35_GBO0;
assign R23C35_GB10 = R23C35_GBO0;
assign R23C36_GB10 = R23C35_GBO0;
assign R23C37_GB10 = R23C35_GBO0;
assign R24C34_GB10 = R24C35_GBO0;
assign R24C35_GB10 = R24C35_GBO0;
assign R24C36_GB10 = R24C35_GBO0;
assign R24C37_GB10 = R24C35_GBO0;
assign R25C34_GB10 = R25C35_GBO0;
assign R25C35_GB10 = R25C35_GBO0;
assign R25C36_GB10 = R25C35_GBO0;
assign R25C37_GB10 = R25C35_GBO0;
assign R26C34_GB10 = R26C35_GBO0;
assign R26C35_GB10 = R26C35_GBO0;
assign R26C36_GB10 = R26C35_GBO0;
assign R26C37_GB10 = R26C35_GBO0;
assign R27C34_GB10 = R27C35_GBO0;
assign R27C35_GB10 = R27C35_GBO0;
assign R27C36_GB10 = R27C35_GBO0;
assign R27C37_GB10 = R27C35_GBO0;
assign R11C41_GB10 = R11C39_GBO0;
assign R11C38_GB10 = R11C39_GBO0;
assign R11C39_GB10 = R11C39_GBO0;
assign R11C40_GB10 = R11C39_GBO0;
assign R12C41_GB10 = R12C39_GBO0;
assign R12C38_GB10 = R12C39_GBO0;
assign R12C39_GB10 = R12C39_GBO0;
assign R12C40_GB10 = R12C39_GBO0;
assign R13C41_GB10 = R13C39_GBO0;
assign R13C38_GB10 = R13C39_GBO0;
assign R13C39_GB10 = R13C39_GBO0;
assign R13C40_GB10 = R13C39_GBO0;
assign R14C41_GB10 = R14C39_GBO0;
assign R14C38_GB10 = R14C39_GBO0;
assign R14C39_GB10 = R14C39_GBO0;
assign R14C40_GB10 = R14C39_GBO0;
assign R15C41_GB10 = R15C39_GBO0;
assign R15C38_GB10 = R15C39_GBO0;
assign R15C39_GB10 = R15C39_GBO0;
assign R15C40_GB10 = R15C39_GBO0;
assign R16C41_GB10 = R16C39_GBO0;
assign R16C38_GB10 = R16C39_GBO0;
assign R16C39_GB10 = R16C39_GBO0;
assign R16C40_GB10 = R16C39_GBO0;
assign R17C41_GB10 = R17C39_GBO0;
assign R17C38_GB10 = R17C39_GBO0;
assign R17C39_GB10 = R17C39_GBO0;
assign R17C40_GB10 = R17C39_GBO0;
assign R18C41_GB10 = R18C39_GBO0;
assign R18C38_GB10 = R18C39_GBO0;
assign R18C39_GB10 = R18C39_GBO0;
assign R18C40_GB10 = R18C39_GBO0;
assign R20C41_GB10 = R20C39_GBO0;
assign R20C38_GB10 = R20C39_GBO0;
assign R20C39_GB10 = R20C39_GBO0;
assign R20C40_GB10 = R20C39_GBO0;
assign R21C41_GB10 = R21C39_GBO0;
assign R21C38_GB10 = R21C39_GBO0;
assign R21C39_GB10 = R21C39_GBO0;
assign R21C40_GB10 = R21C39_GBO0;
assign R22C41_GB10 = R22C39_GBO0;
assign R22C38_GB10 = R22C39_GBO0;
assign R22C39_GB10 = R22C39_GBO0;
assign R22C40_GB10 = R22C39_GBO0;
assign R23C41_GB10 = R23C39_GBO0;
assign R23C38_GB10 = R23C39_GBO0;
assign R23C39_GB10 = R23C39_GBO0;
assign R23C40_GB10 = R23C39_GBO0;
assign R24C41_GB10 = R24C39_GBO0;
assign R24C38_GB10 = R24C39_GBO0;
assign R24C39_GB10 = R24C39_GBO0;
assign R24C40_GB10 = R24C39_GBO0;
assign R25C41_GB10 = R25C39_GBO0;
assign R25C38_GB10 = R25C39_GBO0;
assign R25C39_GB10 = R25C39_GBO0;
assign R25C40_GB10 = R25C39_GBO0;
assign R26C41_GB10 = R26C39_GBO0;
assign R26C38_GB10 = R26C39_GBO0;
assign R26C39_GB10 = R26C39_GBO0;
assign R26C40_GB10 = R26C39_GBO0;
assign R27C41_GB10 = R27C39_GBO0;
assign R27C38_GB10 = R27C39_GBO0;
assign R27C39_GB10 = R27C39_GBO0;
assign R27C40_GB10 = R27C39_GBO0;
assign R11C42_GB10 = R11C43_GBO0;
assign R11C43_GB10 = R11C43_GBO0;
assign R11C44_GB10 = R11C43_GBO0;
assign R11C45_GB10 = R11C43_GBO0;
assign R11C46_GB10 = R11C43_GBO0;
assign R12C42_GB10 = R12C43_GBO0;
assign R12C43_GB10 = R12C43_GBO0;
assign R12C44_GB10 = R12C43_GBO0;
assign R12C45_GB10 = R12C43_GBO0;
assign R12C46_GB10 = R12C43_GBO0;
assign R13C42_GB10 = R13C43_GBO0;
assign R13C43_GB10 = R13C43_GBO0;
assign R13C44_GB10 = R13C43_GBO0;
assign R13C45_GB10 = R13C43_GBO0;
assign R13C46_GB10 = R13C43_GBO0;
assign R14C42_GB10 = R14C43_GBO0;
assign R14C43_GB10 = R14C43_GBO0;
assign R14C44_GB10 = R14C43_GBO0;
assign R14C45_GB10 = R14C43_GBO0;
assign R14C46_GB10 = R14C43_GBO0;
assign R15C42_GB10 = R15C43_GBO0;
assign R15C43_GB10 = R15C43_GBO0;
assign R15C44_GB10 = R15C43_GBO0;
assign R15C45_GB10 = R15C43_GBO0;
assign R15C46_GB10 = R15C43_GBO0;
assign R16C42_GB10 = R16C43_GBO0;
assign R16C43_GB10 = R16C43_GBO0;
assign R16C44_GB10 = R16C43_GBO0;
assign R16C45_GB10 = R16C43_GBO0;
assign R16C46_GB10 = R16C43_GBO0;
assign R17C42_GB10 = R17C43_GBO0;
assign R17C43_GB10 = R17C43_GBO0;
assign R17C44_GB10 = R17C43_GBO0;
assign R17C45_GB10 = R17C43_GBO0;
assign R17C46_GB10 = R17C43_GBO0;
assign R18C42_GB10 = R18C43_GBO0;
assign R18C43_GB10 = R18C43_GBO0;
assign R18C44_GB10 = R18C43_GBO0;
assign R18C45_GB10 = R18C43_GBO0;
assign R18C46_GB10 = R18C43_GBO0;
assign R20C42_GB10 = R20C43_GBO0;
assign R20C43_GB10 = R20C43_GBO0;
assign R20C44_GB10 = R20C43_GBO0;
assign R20C45_GB10 = R20C43_GBO0;
assign R20C46_GB10 = R20C43_GBO0;
assign R21C42_GB10 = R21C43_GBO0;
assign R21C43_GB10 = R21C43_GBO0;
assign R21C44_GB10 = R21C43_GBO0;
assign R21C45_GB10 = R21C43_GBO0;
assign R21C46_GB10 = R21C43_GBO0;
assign R22C42_GB10 = R22C43_GBO0;
assign R22C43_GB10 = R22C43_GBO0;
assign R22C44_GB10 = R22C43_GBO0;
assign R22C45_GB10 = R22C43_GBO0;
assign R22C46_GB10 = R22C43_GBO0;
assign R23C42_GB10 = R23C43_GBO0;
assign R23C43_GB10 = R23C43_GBO0;
assign R23C44_GB10 = R23C43_GBO0;
assign R23C45_GB10 = R23C43_GBO0;
assign R23C46_GB10 = R23C43_GBO0;
assign R24C42_GB10 = R24C43_GBO0;
assign R24C43_GB10 = R24C43_GBO0;
assign R24C44_GB10 = R24C43_GBO0;
assign R24C45_GB10 = R24C43_GBO0;
assign R24C46_GB10 = R24C43_GBO0;
assign R25C42_GB10 = R25C43_GBO0;
assign R25C43_GB10 = R25C43_GBO0;
assign R25C44_GB10 = R25C43_GBO0;
assign R25C45_GB10 = R25C43_GBO0;
assign R25C46_GB10 = R25C43_GBO0;
assign R26C42_GB10 = R26C43_GBO0;
assign R26C43_GB10 = R26C43_GBO0;
assign R26C44_GB10 = R26C43_GBO0;
assign R26C45_GB10 = R26C43_GBO0;
assign R26C46_GB10 = R26C43_GBO0;
assign R27C42_GB10 = R27C43_GBO0;
assign R27C43_GB10 = R27C43_GBO0;
assign R27C44_GB10 = R27C43_GBO0;
assign R27C45_GB10 = R27C43_GBO0;
assign R27C46_GB10 = R27C43_GBO0;
assign R11C29_GB20 = R11C30_GBO0;
assign R11C30_GB20 = R11C30_GBO0;
assign R11C31_GB20 = R11C30_GBO0;
assign R11C32_GB20 = R11C30_GBO0;
assign R12C29_GB20 = R12C30_GBO0;
assign R12C30_GB20 = R12C30_GBO0;
assign R12C31_GB20 = R12C30_GBO0;
assign R12C32_GB20 = R12C30_GBO0;
assign R13C29_GB20 = R13C30_GBO0;
assign R13C30_GB20 = R13C30_GBO0;
assign R13C31_GB20 = R13C30_GBO0;
assign R13C32_GB20 = R13C30_GBO0;
assign R14C29_GB20 = R14C30_GBO0;
assign R14C30_GB20 = R14C30_GBO0;
assign R14C31_GB20 = R14C30_GBO0;
assign R14C32_GB20 = R14C30_GBO0;
assign R15C29_GB20 = R15C30_GBO0;
assign R15C30_GB20 = R15C30_GBO0;
assign R15C31_GB20 = R15C30_GBO0;
assign R15C32_GB20 = R15C30_GBO0;
assign R16C29_GB20 = R16C30_GBO0;
assign R16C30_GB20 = R16C30_GBO0;
assign R16C31_GB20 = R16C30_GBO0;
assign R16C32_GB20 = R16C30_GBO0;
assign R17C29_GB20 = R17C30_GBO0;
assign R17C30_GB20 = R17C30_GBO0;
assign R17C31_GB20 = R17C30_GBO0;
assign R17C32_GB20 = R17C30_GBO0;
assign R18C29_GB20 = R18C30_GBO0;
assign R18C30_GB20 = R18C30_GBO0;
assign R18C31_GB20 = R18C30_GBO0;
assign R18C32_GB20 = R18C30_GBO0;
assign R20C29_GB20 = R20C30_GBO0;
assign R20C30_GB20 = R20C30_GBO0;
assign R20C31_GB20 = R20C30_GBO0;
assign R20C32_GB20 = R20C30_GBO0;
assign R21C29_GB20 = R21C30_GBO0;
assign R21C30_GB20 = R21C30_GBO0;
assign R21C31_GB20 = R21C30_GBO0;
assign R21C32_GB20 = R21C30_GBO0;
assign R22C29_GB20 = R22C30_GBO0;
assign R22C30_GB20 = R22C30_GBO0;
assign R22C31_GB20 = R22C30_GBO0;
assign R22C32_GB20 = R22C30_GBO0;
assign R23C29_GB20 = R23C30_GBO0;
assign R23C30_GB20 = R23C30_GBO0;
assign R23C31_GB20 = R23C30_GBO0;
assign R23C32_GB20 = R23C30_GBO0;
assign R24C29_GB20 = R24C30_GBO0;
assign R24C30_GB20 = R24C30_GBO0;
assign R24C31_GB20 = R24C30_GBO0;
assign R24C32_GB20 = R24C30_GBO0;
assign R25C29_GB20 = R25C30_GBO0;
assign R25C30_GB20 = R25C30_GBO0;
assign R25C31_GB20 = R25C30_GBO0;
assign R25C32_GB20 = R25C30_GBO0;
assign R26C29_GB20 = R26C30_GBO0;
assign R26C30_GB20 = R26C30_GBO0;
assign R26C31_GB20 = R26C30_GBO0;
assign R26C32_GB20 = R26C30_GBO0;
assign R27C29_GB20 = R27C30_GBO0;
assign R27C30_GB20 = R27C30_GBO0;
assign R27C31_GB20 = R27C30_GBO0;
assign R27C32_GB20 = R27C30_GBO0;
assign R11C33_GB20 = R11C34_GBO0;
assign R11C34_GB20 = R11C34_GBO0;
assign R11C35_GB20 = R11C34_GBO0;
assign R11C36_GB20 = R11C34_GBO0;
assign R12C33_GB20 = R12C34_GBO0;
assign R12C34_GB20 = R12C34_GBO0;
assign R12C35_GB20 = R12C34_GBO0;
assign R12C36_GB20 = R12C34_GBO0;
assign R13C33_GB20 = R13C34_GBO0;
assign R13C34_GB20 = R13C34_GBO0;
assign R13C35_GB20 = R13C34_GBO0;
assign R13C36_GB20 = R13C34_GBO0;
assign R14C33_GB20 = R14C34_GBO0;
assign R14C34_GB20 = R14C34_GBO0;
assign R14C35_GB20 = R14C34_GBO0;
assign R14C36_GB20 = R14C34_GBO0;
assign R15C33_GB20 = R15C34_GBO0;
assign R15C34_GB20 = R15C34_GBO0;
assign R15C35_GB20 = R15C34_GBO0;
assign R15C36_GB20 = R15C34_GBO0;
assign R16C33_GB20 = R16C34_GBO0;
assign R16C34_GB20 = R16C34_GBO0;
assign R16C35_GB20 = R16C34_GBO0;
assign R16C36_GB20 = R16C34_GBO0;
assign R17C33_GB20 = R17C34_GBO0;
assign R17C34_GB20 = R17C34_GBO0;
assign R17C35_GB20 = R17C34_GBO0;
assign R17C36_GB20 = R17C34_GBO0;
assign R18C33_GB20 = R18C34_GBO0;
assign R18C34_GB20 = R18C34_GBO0;
assign R18C35_GB20 = R18C34_GBO0;
assign R18C36_GB20 = R18C34_GBO0;
assign R20C33_GB20 = R20C34_GBO0;
assign R20C34_GB20 = R20C34_GBO0;
assign R20C35_GB20 = R20C34_GBO0;
assign R20C36_GB20 = R20C34_GBO0;
assign R21C33_GB20 = R21C34_GBO0;
assign R21C34_GB20 = R21C34_GBO0;
assign R21C35_GB20 = R21C34_GBO0;
assign R21C36_GB20 = R21C34_GBO0;
assign R22C33_GB20 = R22C34_GBO0;
assign R22C34_GB20 = R22C34_GBO0;
assign R22C35_GB20 = R22C34_GBO0;
assign R22C36_GB20 = R22C34_GBO0;
assign R23C33_GB20 = R23C34_GBO0;
assign R23C34_GB20 = R23C34_GBO0;
assign R23C35_GB20 = R23C34_GBO0;
assign R23C36_GB20 = R23C34_GBO0;
assign R24C33_GB20 = R24C34_GBO0;
assign R24C34_GB20 = R24C34_GBO0;
assign R24C35_GB20 = R24C34_GBO0;
assign R24C36_GB20 = R24C34_GBO0;
assign R25C33_GB20 = R25C34_GBO0;
assign R25C34_GB20 = R25C34_GBO0;
assign R25C35_GB20 = R25C34_GBO0;
assign R25C36_GB20 = R25C34_GBO0;
assign R26C33_GB20 = R26C34_GBO0;
assign R26C34_GB20 = R26C34_GBO0;
assign R26C35_GB20 = R26C34_GBO0;
assign R26C36_GB20 = R26C34_GBO0;
assign R27C33_GB20 = R27C34_GBO0;
assign R27C34_GB20 = R27C34_GBO0;
assign R27C35_GB20 = R27C34_GBO0;
assign R27C36_GB20 = R27C34_GBO0;
assign R11C37_GB20 = R11C38_GBO0;
assign R11C38_GB20 = R11C38_GBO0;
assign R11C39_GB20 = R11C38_GBO0;
assign R11C40_GB20 = R11C38_GBO0;
assign R12C37_GB20 = R12C38_GBO0;
assign R12C38_GB20 = R12C38_GBO0;
assign R12C39_GB20 = R12C38_GBO0;
assign R12C40_GB20 = R12C38_GBO0;
assign R13C37_GB20 = R13C38_GBO0;
assign R13C38_GB20 = R13C38_GBO0;
assign R13C39_GB20 = R13C38_GBO0;
assign R13C40_GB20 = R13C38_GBO0;
assign R14C37_GB20 = R14C38_GBO0;
assign R14C38_GB20 = R14C38_GBO0;
assign R14C39_GB20 = R14C38_GBO0;
assign R14C40_GB20 = R14C38_GBO0;
assign R15C37_GB20 = R15C38_GBO0;
assign R15C38_GB20 = R15C38_GBO0;
assign R15C39_GB20 = R15C38_GBO0;
assign R15C40_GB20 = R15C38_GBO0;
assign R16C37_GB20 = R16C38_GBO0;
assign R16C38_GB20 = R16C38_GBO0;
assign R16C39_GB20 = R16C38_GBO0;
assign R16C40_GB20 = R16C38_GBO0;
assign R17C37_GB20 = R17C38_GBO0;
assign R17C38_GB20 = R17C38_GBO0;
assign R17C39_GB20 = R17C38_GBO0;
assign R17C40_GB20 = R17C38_GBO0;
assign R18C37_GB20 = R18C38_GBO0;
assign R18C38_GB20 = R18C38_GBO0;
assign R18C39_GB20 = R18C38_GBO0;
assign R18C40_GB20 = R18C38_GBO0;
assign R20C37_GB20 = R20C38_GBO0;
assign R20C38_GB20 = R20C38_GBO0;
assign R20C39_GB20 = R20C38_GBO0;
assign R20C40_GB20 = R20C38_GBO0;
assign R21C37_GB20 = R21C38_GBO0;
assign R21C38_GB20 = R21C38_GBO0;
assign R21C39_GB20 = R21C38_GBO0;
assign R21C40_GB20 = R21C38_GBO0;
assign R22C37_GB20 = R22C38_GBO0;
assign R22C38_GB20 = R22C38_GBO0;
assign R22C39_GB20 = R22C38_GBO0;
assign R22C40_GB20 = R22C38_GBO0;
assign R23C37_GB20 = R23C38_GBO0;
assign R23C38_GB20 = R23C38_GBO0;
assign R23C39_GB20 = R23C38_GBO0;
assign R23C40_GB20 = R23C38_GBO0;
assign R24C37_GB20 = R24C38_GBO0;
assign R24C38_GB20 = R24C38_GBO0;
assign R24C39_GB20 = R24C38_GBO0;
assign R24C40_GB20 = R24C38_GBO0;
assign R25C37_GB20 = R25C38_GBO0;
assign R25C38_GB20 = R25C38_GBO0;
assign R25C39_GB20 = R25C38_GBO0;
assign R25C40_GB20 = R25C38_GBO0;
assign R26C37_GB20 = R26C38_GBO0;
assign R26C38_GB20 = R26C38_GBO0;
assign R26C39_GB20 = R26C38_GBO0;
assign R26C40_GB20 = R26C38_GBO0;
assign R27C37_GB20 = R27C38_GBO0;
assign R27C38_GB20 = R27C38_GBO0;
assign R27C39_GB20 = R27C38_GBO0;
assign R27C40_GB20 = R27C38_GBO0;
assign R11C41_GB20 = R11C42_GBO0;
assign R11C42_GB20 = R11C42_GBO0;
assign R11C43_GB20 = R11C42_GBO0;
assign R11C44_GB20 = R11C42_GBO0;
assign R12C41_GB20 = R12C42_GBO0;
assign R12C42_GB20 = R12C42_GBO0;
assign R12C43_GB20 = R12C42_GBO0;
assign R12C44_GB20 = R12C42_GBO0;
assign R13C41_GB20 = R13C42_GBO0;
assign R13C42_GB20 = R13C42_GBO0;
assign R13C43_GB20 = R13C42_GBO0;
assign R13C44_GB20 = R13C42_GBO0;
assign R14C41_GB20 = R14C42_GBO0;
assign R14C42_GB20 = R14C42_GBO0;
assign R14C43_GB20 = R14C42_GBO0;
assign R14C44_GB20 = R14C42_GBO0;
assign R15C41_GB20 = R15C42_GBO0;
assign R15C42_GB20 = R15C42_GBO0;
assign R15C43_GB20 = R15C42_GBO0;
assign R15C44_GB20 = R15C42_GBO0;
assign R16C41_GB20 = R16C42_GBO0;
assign R16C42_GB20 = R16C42_GBO0;
assign R16C43_GB20 = R16C42_GBO0;
assign R16C44_GB20 = R16C42_GBO0;
assign R17C41_GB20 = R17C42_GBO0;
assign R17C42_GB20 = R17C42_GBO0;
assign R17C43_GB20 = R17C42_GBO0;
assign R17C44_GB20 = R17C42_GBO0;
assign R18C41_GB20 = R18C42_GBO0;
assign R18C42_GB20 = R18C42_GBO0;
assign R18C43_GB20 = R18C42_GBO0;
assign R18C44_GB20 = R18C42_GBO0;
assign R20C41_GB20 = R20C42_GBO0;
assign R20C42_GB20 = R20C42_GBO0;
assign R20C43_GB20 = R20C42_GBO0;
assign R20C44_GB20 = R20C42_GBO0;
assign R21C41_GB20 = R21C42_GBO0;
assign R21C42_GB20 = R21C42_GBO0;
assign R21C43_GB20 = R21C42_GBO0;
assign R21C44_GB20 = R21C42_GBO0;
assign R22C41_GB20 = R22C42_GBO0;
assign R22C42_GB20 = R22C42_GBO0;
assign R22C43_GB20 = R22C42_GBO0;
assign R22C44_GB20 = R22C42_GBO0;
assign R23C41_GB20 = R23C42_GBO0;
assign R23C42_GB20 = R23C42_GBO0;
assign R23C43_GB20 = R23C42_GBO0;
assign R23C44_GB20 = R23C42_GBO0;
assign R24C41_GB20 = R24C42_GBO0;
assign R24C42_GB20 = R24C42_GBO0;
assign R24C43_GB20 = R24C42_GBO0;
assign R24C44_GB20 = R24C42_GBO0;
assign R25C41_GB20 = R25C42_GBO0;
assign R25C42_GB20 = R25C42_GBO0;
assign R25C43_GB20 = R25C42_GBO0;
assign R25C44_GB20 = R25C42_GBO0;
assign R26C41_GB20 = R26C42_GBO0;
assign R26C42_GB20 = R26C42_GBO0;
assign R26C43_GB20 = R26C42_GBO0;
assign R26C44_GB20 = R26C42_GBO0;
assign R27C41_GB20 = R27C42_GBO0;
assign R27C42_GB20 = R27C42_GBO0;
assign R27C43_GB20 = R27C42_GBO0;
assign R27C44_GB20 = R27C42_GBO0;
assign R11C45_GB20 = R11C46_GBO0;
assign R11C46_GB20 = R11C46_GBO0;
assign R12C45_GB20 = R12C46_GBO0;
assign R12C46_GB20 = R12C46_GBO0;
assign R13C45_GB20 = R13C46_GBO0;
assign R13C46_GB20 = R13C46_GBO0;
assign R14C45_GB20 = R14C46_GBO0;
assign R14C46_GB20 = R14C46_GBO0;
assign R15C45_GB20 = R15C46_GBO0;
assign R15C46_GB20 = R15C46_GBO0;
assign R16C45_GB20 = R16C46_GBO0;
assign R16C46_GB20 = R16C46_GBO0;
assign R17C45_GB20 = R17C46_GBO0;
assign R17C46_GB20 = R17C46_GBO0;
assign R18C45_GB20 = R18C46_GBO0;
assign R18C46_GB20 = R18C46_GBO0;
assign R20C45_GB20 = R20C46_GBO0;
assign R20C46_GB20 = R20C46_GBO0;
assign R21C45_GB20 = R21C46_GBO0;
assign R21C46_GB20 = R21C46_GBO0;
assign R22C45_GB20 = R22C46_GBO0;
assign R22C46_GB20 = R22C46_GBO0;
assign R23C45_GB20 = R23C46_GBO0;
assign R23C46_GB20 = R23C46_GBO0;
assign R24C45_GB20 = R24C46_GBO0;
assign R24C46_GB20 = R24C46_GBO0;
assign R25C45_GB20 = R25C46_GBO0;
assign R25C46_GB20 = R25C46_GBO0;
assign R26C45_GB20 = R26C46_GBO0;
assign R26C46_GB20 = R26C46_GBO0;
assign R27C45_GB20 = R27C46_GBO0;
assign R27C46_GB20 = R27C46_GBO0;
assign R11C29_GB30 = R11C29_GBO0;
assign R11C30_GB30 = R11C29_GBO0;
assign R11C31_GB30 = R11C29_GBO0;
assign R12C29_GB30 = R12C29_GBO0;
assign R12C30_GB30 = R12C29_GBO0;
assign R12C31_GB30 = R12C29_GBO0;
assign R13C29_GB30 = R13C29_GBO0;
assign R13C30_GB30 = R13C29_GBO0;
assign R13C31_GB30 = R13C29_GBO0;
assign R14C29_GB30 = R14C29_GBO0;
assign R14C30_GB30 = R14C29_GBO0;
assign R14C31_GB30 = R14C29_GBO0;
assign R15C29_GB30 = R15C29_GBO0;
assign R15C30_GB30 = R15C29_GBO0;
assign R15C31_GB30 = R15C29_GBO0;
assign R16C29_GB30 = R16C29_GBO0;
assign R16C30_GB30 = R16C29_GBO0;
assign R16C31_GB30 = R16C29_GBO0;
assign R17C29_GB30 = R17C29_GBO0;
assign R17C30_GB30 = R17C29_GBO0;
assign R17C31_GB30 = R17C29_GBO0;
assign R18C29_GB30 = R18C29_GBO0;
assign R18C30_GB30 = R18C29_GBO0;
assign R18C31_GB30 = R18C29_GBO0;
assign R20C29_GB30 = R20C29_GBO0;
assign R20C30_GB30 = R20C29_GBO0;
assign R20C31_GB30 = R20C29_GBO0;
assign R21C29_GB30 = R21C29_GBO0;
assign R21C30_GB30 = R21C29_GBO0;
assign R21C31_GB30 = R21C29_GBO0;
assign R22C29_GB30 = R22C29_GBO0;
assign R22C30_GB30 = R22C29_GBO0;
assign R22C31_GB30 = R22C29_GBO0;
assign R23C29_GB30 = R23C29_GBO0;
assign R23C30_GB30 = R23C29_GBO0;
assign R23C31_GB30 = R23C29_GBO0;
assign R24C29_GB30 = R24C29_GBO0;
assign R24C30_GB30 = R24C29_GBO0;
assign R24C31_GB30 = R24C29_GBO0;
assign R25C29_GB30 = R25C29_GBO0;
assign R25C30_GB30 = R25C29_GBO0;
assign R25C31_GB30 = R25C29_GBO0;
assign R26C29_GB30 = R26C29_GBO0;
assign R26C30_GB30 = R26C29_GBO0;
assign R26C31_GB30 = R26C29_GBO0;
assign R27C29_GB30 = R27C29_GBO0;
assign R27C30_GB30 = R27C29_GBO0;
assign R27C31_GB30 = R27C29_GBO0;
assign R11C33_GB30 = R11C33_GBO0;
assign R11C34_GB30 = R11C33_GBO0;
assign R11C35_GB30 = R11C33_GBO0;
assign R11C32_GB30 = R11C33_GBO0;
assign R12C33_GB30 = R12C33_GBO0;
assign R12C34_GB30 = R12C33_GBO0;
assign R12C35_GB30 = R12C33_GBO0;
assign R12C32_GB30 = R12C33_GBO0;
assign R13C33_GB30 = R13C33_GBO0;
assign R13C34_GB30 = R13C33_GBO0;
assign R13C35_GB30 = R13C33_GBO0;
assign R13C32_GB30 = R13C33_GBO0;
assign R14C33_GB30 = R14C33_GBO0;
assign R14C34_GB30 = R14C33_GBO0;
assign R14C35_GB30 = R14C33_GBO0;
assign R14C32_GB30 = R14C33_GBO0;
assign R15C33_GB30 = R15C33_GBO0;
assign R15C34_GB30 = R15C33_GBO0;
assign R15C35_GB30 = R15C33_GBO0;
assign R15C32_GB30 = R15C33_GBO0;
assign R16C33_GB30 = R16C33_GBO0;
assign R16C34_GB30 = R16C33_GBO0;
assign R16C35_GB30 = R16C33_GBO0;
assign R16C32_GB30 = R16C33_GBO0;
assign R17C33_GB30 = R17C33_GBO0;
assign R17C34_GB30 = R17C33_GBO0;
assign R17C35_GB30 = R17C33_GBO0;
assign R17C32_GB30 = R17C33_GBO0;
assign R18C33_GB30 = R18C33_GBO0;
assign R18C34_GB30 = R18C33_GBO0;
assign R18C35_GB30 = R18C33_GBO0;
assign R18C32_GB30 = R18C33_GBO0;
assign R20C33_GB30 = R20C33_GBO0;
assign R20C34_GB30 = R20C33_GBO0;
assign R20C35_GB30 = R20C33_GBO0;
assign R20C32_GB30 = R20C33_GBO0;
assign R21C33_GB30 = R21C33_GBO0;
assign R21C34_GB30 = R21C33_GBO0;
assign R21C35_GB30 = R21C33_GBO0;
assign R21C32_GB30 = R21C33_GBO0;
assign R22C33_GB30 = R22C33_GBO0;
assign R22C34_GB30 = R22C33_GBO0;
assign R22C35_GB30 = R22C33_GBO0;
assign R22C32_GB30 = R22C33_GBO0;
assign R23C33_GB30 = R23C33_GBO0;
assign R23C34_GB30 = R23C33_GBO0;
assign R23C35_GB30 = R23C33_GBO0;
assign R23C32_GB30 = R23C33_GBO0;
assign R24C33_GB30 = R24C33_GBO0;
assign R24C34_GB30 = R24C33_GBO0;
assign R24C35_GB30 = R24C33_GBO0;
assign R24C32_GB30 = R24C33_GBO0;
assign R25C33_GB30 = R25C33_GBO0;
assign R25C34_GB30 = R25C33_GBO0;
assign R25C35_GB30 = R25C33_GBO0;
assign R25C32_GB30 = R25C33_GBO0;
assign R26C33_GB30 = R26C33_GBO0;
assign R26C34_GB30 = R26C33_GBO0;
assign R26C35_GB30 = R26C33_GBO0;
assign R26C32_GB30 = R26C33_GBO0;
assign R27C33_GB30 = R27C33_GBO0;
assign R27C34_GB30 = R27C33_GBO0;
assign R27C35_GB30 = R27C33_GBO0;
assign R27C32_GB30 = R27C33_GBO0;
assign R11C36_GB30 = R11C37_GBO0;
assign R11C37_GB30 = R11C37_GBO0;
assign R11C38_GB30 = R11C37_GBO0;
assign R11C39_GB30 = R11C37_GBO0;
assign R12C36_GB30 = R12C37_GBO0;
assign R12C37_GB30 = R12C37_GBO0;
assign R12C38_GB30 = R12C37_GBO0;
assign R12C39_GB30 = R12C37_GBO0;
assign R13C36_GB30 = R13C37_GBO0;
assign R13C37_GB30 = R13C37_GBO0;
assign R13C38_GB30 = R13C37_GBO0;
assign R13C39_GB30 = R13C37_GBO0;
assign R14C36_GB30 = R14C37_GBO0;
assign R14C37_GB30 = R14C37_GBO0;
assign R14C38_GB30 = R14C37_GBO0;
assign R14C39_GB30 = R14C37_GBO0;
assign R15C36_GB30 = R15C37_GBO0;
assign R15C37_GB30 = R15C37_GBO0;
assign R15C38_GB30 = R15C37_GBO0;
assign R15C39_GB30 = R15C37_GBO0;
assign R16C36_GB30 = R16C37_GBO0;
assign R16C37_GB30 = R16C37_GBO0;
assign R16C38_GB30 = R16C37_GBO0;
assign R16C39_GB30 = R16C37_GBO0;
assign R17C36_GB30 = R17C37_GBO0;
assign R17C37_GB30 = R17C37_GBO0;
assign R17C38_GB30 = R17C37_GBO0;
assign R17C39_GB30 = R17C37_GBO0;
assign R18C36_GB30 = R18C37_GBO0;
assign R18C37_GB30 = R18C37_GBO0;
assign R18C38_GB30 = R18C37_GBO0;
assign R18C39_GB30 = R18C37_GBO0;
assign R20C36_GB30 = R20C37_GBO0;
assign R20C37_GB30 = R20C37_GBO0;
assign R20C38_GB30 = R20C37_GBO0;
assign R20C39_GB30 = R20C37_GBO0;
assign R21C36_GB30 = R21C37_GBO0;
assign R21C37_GB30 = R21C37_GBO0;
assign R21C38_GB30 = R21C37_GBO0;
assign R21C39_GB30 = R21C37_GBO0;
assign R22C36_GB30 = R22C37_GBO0;
assign R22C37_GB30 = R22C37_GBO0;
assign R22C38_GB30 = R22C37_GBO0;
assign R22C39_GB30 = R22C37_GBO0;
assign R23C36_GB30 = R23C37_GBO0;
assign R23C37_GB30 = R23C37_GBO0;
assign R23C38_GB30 = R23C37_GBO0;
assign R23C39_GB30 = R23C37_GBO0;
assign R24C36_GB30 = R24C37_GBO0;
assign R24C37_GB30 = R24C37_GBO0;
assign R24C38_GB30 = R24C37_GBO0;
assign R24C39_GB30 = R24C37_GBO0;
assign R25C36_GB30 = R25C37_GBO0;
assign R25C37_GB30 = R25C37_GBO0;
assign R25C38_GB30 = R25C37_GBO0;
assign R25C39_GB30 = R25C37_GBO0;
assign R26C36_GB30 = R26C37_GBO0;
assign R26C37_GB30 = R26C37_GBO0;
assign R26C38_GB30 = R26C37_GBO0;
assign R26C39_GB30 = R26C37_GBO0;
assign R27C36_GB30 = R27C37_GBO0;
assign R27C37_GB30 = R27C37_GBO0;
assign R27C38_GB30 = R27C37_GBO0;
assign R27C39_GB30 = R27C37_GBO0;
assign R11C41_GB30 = R11C41_GBO0;
assign R11C42_GB30 = R11C41_GBO0;
assign R11C43_GB30 = R11C41_GBO0;
assign R11C40_GB30 = R11C41_GBO0;
assign R12C41_GB30 = R12C41_GBO0;
assign R12C42_GB30 = R12C41_GBO0;
assign R12C43_GB30 = R12C41_GBO0;
assign R12C40_GB30 = R12C41_GBO0;
assign R13C41_GB30 = R13C41_GBO0;
assign R13C42_GB30 = R13C41_GBO0;
assign R13C43_GB30 = R13C41_GBO0;
assign R13C40_GB30 = R13C41_GBO0;
assign R14C41_GB30 = R14C41_GBO0;
assign R14C42_GB30 = R14C41_GBO0;
assign R14C43_GB30 = R14C41_GBO0;
assign R14C40_GB30 = R14C41_GBO0;
assign R15C41_GB30 = R15C41_GBO0;
assign R15C42_GB30 = R15C41_GBO0;
assign R15C43_GB30 = R15C41_GBO0;
assign R15C40_GB30 = R15C41_GBO0;
assign R16C41_GB30 = R16C41_GBO0;
assign R16C42_GB30 = R16C41_GBO0;
assign R16C43_GB30 = R16C41_GBO0;
assign R16C40_GB30 = R16C41_GBO0;
assign R17C41_GB30 = R17C41_GBO0;
assign R17C42_GB30 = R17C41_GBO0;
assign R17C43_GB30 = R17C41_GBO0;
assign R17C40_GB30 = R17C41_GBO0;
assign R18C41_GB30 = R18C41_GBO0;
assign R18C42_GB30 = R18C41_GBO0;
assign R18C43_GB30 = R18C41_GBO0;
assign R18C40_GB30 = R18C41_GBO0;
assign R20C41_GB30 = R20C41_GBO0;
assign R20C42_GB30 = R20C41_GBO0;
assign R20C43_GB30 = R20C41_GBO0;
assign R20C40_GB30 = R20C41_GBO0;
assign R21C41_GB30 = R21C41_GBO0;
assign R21C42_GB30 = R21C41_GBO0;
assign R21C43_GB30 = R21C41_GBO0;
assign R21C40_GB30 = R21C41_GBO0;
assign R22C41_GB30 = R22C41_GBO0;
assign R22C42_GB30 = R22C41_GBO0;
assign R22C43_GB30 = R22C41_GBO0;
assign R22C40_GB30 = R22C41_GBO0;
assign R23C41_GB30 = R23C41_GBO0;
assign R23C42_GB30 = R23C41_GBO0;
assign R23C43_GB30 = R23C41_GBO0;
assign R23C40_GB30 = R23C41_GBO0;
assign R24C41_GB30 = R24C41_GBO0;
assign R24C42_GB30 = R24C41_GBO0;
assign R24C43_GB30 = R24C41_GBO0;
assign R24C40_GB30 = R24C41_GBO0;
assign R25C41_GB30 = R25C41_GBO0;
assign R25C42_GB30 = R25C41_GBO0;
assign R25C43_GB30 = R25C41_GBO0;
assign R25C40_GB30 = R25C41_GBO0;
assign R26C41_GB30 = R26C41_GBO0;
assign R26C42_GB30 = R26C41_GBO0;
assign R26C43_GB30 = R26C41_GBO0;
assign R26C40_GB30 = R26C41_GBO0;
assign R27C41_GB30 = R27C41_GBO0;
assign R27C42_GB30 = R27C41_GBO0;
assign R27C43_GB30 = R27C41_GBO0;
assign R27C40_GB30 = R27C41_GBO0;
assign R11C44_GB30 = R11C45_GBO0;
assign R11C45_GB30 = R11C45_GBO0;
assign R11C46_GB30 = R11C45_GBO0;
assign R12C44_GB30 = R12C45_GBO0;
assign R12C45_GB30 = R12C45_GBO0;
assign R12C46_GB30 = R12C45_GBO0;
assign R13C44_GB30 = R13C45_GBO0;
assign R13C45_GB30 = R13C45_GBO0;
assign R13C46_GB30 = R13C45_GBO0;
assign R14C44_GB30 = R14C45_GBO0;
assign R14C45_GB30 = R14C45_GBO0;
assign R14C46_GB30 = R14C45_GBO0;
assign R15C44_GB30 = R15C45_GBO0;
assign R15C45_GB30 = R15C45_GBO0;
assign R15C46_GB30 = R15C45_GBO0;
assign R16C44_GB30 = R16C45_GBO0;
assign R16C45_GB30 = R16C45_GBO0;
assign R16C46_GB30 = R16C45_GBO0;
assign R17C44_GB30 = R17C45_GBO0;
assign R17C45_GB30 = R17C45_GBO0;
assign R17C46_GB30 = R17C45_GBO0;
assign R18C44_GB30 = R18C45_GBO0;
assign R18C45_GB30 = R18C45_GBO0;
assign R18C46_GB30 = R18C45_GBO0;
assign R20C44_GB30 = R20C45_GBO0;
assign R20C45_GB30 = R20C45_GBO0;
assign R20C46_GB30 = R20C45_GBO0;
assign R21C44_GB30 = R21C45_GBO0;
assign R21C45_GB30 = R21C45_GBO0;
assign R21C46_GB30 = R21C45_GBO0;
assign R22C44_GB30 = R22C45_GBO0;
assign R22C45_GB30 = R22C45_GBO0;
assign R22C46_GB30 = R22C45_GBO0;
assign R23C44_GB30 = R23C45_GBO0;
assign R23C45_GB30 = R23C45_GBO0;
assign R23C46_GB30 = R23C45_GBO0;
assign R24C44_GB30 = R24C45_GBO0;
assign R24C45_GB30 = R24C45_GBO0;
assign R24C46_GB30 = R24C45_GBO0;
assign R25C44_GB30 = R25C45_GBO0;
assign R25C45_GB30 = R25C45_GBO0;
assign R25C46_GB30 = R25C45_GBO0;
assign R26C44_GB30 = R26C45_GBO0;
assign R26C45_GB30 = R26C45_GBO0;
assign R26C46_GB30 = R26C45_GBO0;
assign R27C44_GB30 = R27C45_GBO0;
assign R27C45_GB30 = R27C45_GBO0;
assign R27C46_GB30 = R27C45_GBO0;
assign R11C33_GB40 = R11C32_GBO1;
assign R11C34_GB40 = R11C32_GBO1;
assign R11C29_GB40 = R11C32_GBO1;
assign R11C30_GB40 = R11C32_GBO1;
assign R11C31_GB40 = R11C32_GBO1;
assign R11C32_GB40 = R11C32_GBO1;
assign R12C33_GB40 = R12C32_GBO1;
assign R12C34_GB40 = R12C32_GBO1;
assign R12C29_GB40 = R12C32_GBO1;
assign R12C30_GB40 = R12C32_GBO1;
assign R12C31_GB40 = R12C32_GBO1;
assign R12C32_GB40 = R12C32_GBO1;
assign R13C33_GB40 = R13C32_GBO1;
assign R13C34_GB40 = R13C32_GBO1;
assign R13C29_GB40 = R13C32_GBO1;
assign R13C30_GB40 = R13C32_GBO1;
assign R13C31_GB40 = R13C32_GBO1;
assign R13C32_GB40 = R13C32_GBO1;
assign R14C33_GB40 = R14C32_GBO1;
assign R14C34_GB40 = R14C32_GBO1;
assign R14C29_GB40 = R14C32_GBO1;
assign R14C30_GB40 = R14C32_GBO1;
assign R14C31_GB40 = R14C32_GBO1;
assign R14C32_GB40 = R14C32_GBO1;
assign R15C33_GB40 = R15C32_GBO1;
assign R15C34_GB40 = R15C32_GBO1;
assign R15C29_GB40 = R15C32_GBO1;
assign R15C30_GB40 = R15C32_GBO1;
assign R15C31_GB40 = R15C32_GBO1;
assign R15C32_GB40 = R15C32_GBO1;
assign R16C33_GB40 = R16C32_GBO1;
assign R16C34_GB40 = R16C32_GBO1;
assign R16C29_GB40 = R16C32_GBO1;
assign R16C30_GB40 = R16C32_GBO1;
assign R16C31_GB40 = R16C32_GBO1;
assign R16C32_GB40 = R16C32_GBO1;
assign R17C33_GB40 = R17C32_GBO1;
assign R17C34_GB40 = R17C32_GBO1;
assign R17C29_GB40 = R17C32_GBO1;
assign R17C30_GB40 = R17C32_GBO1;
assign R17C31_GB40 = R17C32_GBO1;
assign R17C32_GB40 = R17C32_GBO1;
assign R18C33_GB40 = R18C32_GBO1;
assign R18C34_GB40 = R18C32_GBO1;
assign R18C29_GB40 = R18C32_GBO1;
assign R18C30_GB40 = R18C32_GBO1;
assign R18C31_GB40 = R18C32_GBO1;
assign R18C32_GB40 = R18C32_GBO1;
assign R20C33_GB40 = R20C32_GBO1;
assign R20C34_GB40 = R20C32_GBO1;
assign R20C29_GB40 = R20C32_GBO1;
assign R20C30_GB40 = R20C32_GBO1;
assign R20C31_GB40 = R20C32_GBO1;
assign R20C32_GB40 = R20C32_GBO1;
assign R21C33_GB40 = R21C32_GBO1;
assign R21C34_GB40 = R21C32_GBO1;
assign R21C29_GB40 = R21C32_GBO1;
assign R21C30_GB40 = R21C32_GBO1;
assign R21C31_GB40 = R21C32_GBO1;
assign R21C32_GB40 = R21C32_GBO1;
assign R22C33_GB40 = R22C32_GBO1;
assign R22C34_GB40 = R22C32_GBO1;
assign R22C29_GB40 = R22C32_GBO1;
assign R22C30_GB40 = R22C32_GBO1;
assign R22C31_GB40 = R22C32_GBO1;
assign R22C32_GB40 = R22C32_GBO1;
assign R23C33_GB40 = R23C32_GBO1;
assign R23C34_GB40 = R23C32_GBO1;
assign R23C29_GB40 = R23C32_GBO1;
assign R23C30_GB40 = R23C32_GBO1;
assign R23C31_GB40 = R23C32_GBO1;
assign R23C32_GB40 = R23C32_GBO1;
assign R24C33_GB40 = R24C32_GBO1;
assign R24C34_GB40 = R24C32_GBO1;
assign R24C29_GB40 = R24C32_GBO1;
assign R24C30_GB40 = R24C32_GBO1;
assign R24C31_GB40 = R24C32_GBO1;
assign R24C32_GB40 = R24C32_GBO1;
assign R25C33_GB40 = R25C32_GBO1;
assign R25C34_GB40 = R25C32_GBO1;
assign R25C29_GB40 = R25C32_GBO1;
assign R25C30_GB40 = R25C32_GBO1;
assign R25C31_GB40 = R25C32_GBO1;
assign R25C32_GB40 = R25C32_GBO1;
assign R26C33_GB40 = R26C32_GBO1;
assign R26C34_GB40 = R26C32_GBO1;
assign R26C29_GB40 = R26C32_GBO1;
assign R26C30_GB40 = R26C32_GBO1;
assign R26C31_GB40 = R26C32_GBO1;
assign R26C32_GB40 = R26C32_GBO1;
assign R27C33_GB40 = R27C32_GBO1;
assign R27C34_GB40 = R27C32_GBO1;
assign R27C29_GB40 = R27C32_GBO1;
assign R27C30_GB40 = R27C32_GBO1;
assign R27C31_GB40 = R27C32_GBO1;
assign R27C32_GB40 = R27C32_GBO1;
assign R11C35_GB40 = R11C36_GBO1;
assign R11C36_GB40 = R11C36_GBO1;
assign R11C37_GB40 = R11C36_GBO1;
assign R11C38_GB40 = R11C36_GBO1;
assign R12C35_GB40 = R12C36_GBO1;
assign R12C36_GB40 = R12C36_GBO1;
assign R12C37_GB40 = R12C36_GBO1;
assign R12C38_GB40 = R12C36_GBO1;
assign R13C35_GB40 = R13C36_GBO1;
assign R13C36_GB40 = R13C36_GBO1;
assign R13C37_GB40 = R13C36_GBO1;
assign R13C38_GB40 = R13C36_GBO1;
assign R14C35_GB40 = R14C36_GBO1;
assign R14C36_GB40 = R14C36_GBO1;
assign R14C37_GB40 = R14C36_GBO1;
assign R14C38_GB40 = R14C36_GBO1;
assign R15C35_GB40 = R15C36_GBO1;
assign R15C36_GB40 = R15C36_GBO1;
assign R15C37_GB40 = R15C36_GBO1;
assign R15C38_GB40 = R15C36_GBO1;
assign R16C35_GB40 = R16C36_GBO1;
assign R16C36_GB40 = R16C36_GBO1;
assign R16C37_GB40 = R16C36_GBO1;
assign R16C38_GB40 = R16C36_GBO1;
assign R17C35_GB40 = R17C36_GBO1;
assign R17C36_GB40 = R17C36_GBO1;
assign R17C37_GB40 = R17C36_GBO1;
assign R17C38_GB40 = R17C36_GBO1;
assign R18C35_GB40 = R18C36_GBO1;
assign R18C36_GB40 = R18C36_GBO1;
assign R18C37_GB40 = R18C36_GBO1;
assign R18C38_GB40 = R18C36_GBO1;
assign R20C35_GB40 = R20C36_GBO1;
assign R20C36_GB40 = R20C36_GBO1;
assign R20C37_GB40 = R20C36_GBO1;
assign R20C38_GB40 = R20C36_GBO1;
assign R21C35_GB40 = R21C36_GBO1;
assign R21C36_GB40 = R21C36_GBO1;
assign R21C37_GB40 = R21C36_GBO1;
assign R21C38_GB40 = R21C36_GBO1;
assign R22C35_GB40 = R22C36_GBO1;
assign R22C36_GB40 = R22C36_GBO1;
assign R22C37_GB40 = R22C36_GBO1;
assign R22C38_GB40 = R22C36_GBO1;
assign R23C35_GB40 = R23C36_GBO1;
assign R23C36_GB40 = R23C36_GBO1;
assign R23C37_GB40 = R23C36_GBO1;
assign R23C38_GB40 = R23C36_GBO1;
assign R24C35_GB40 = R24C36_GBO1;
assign R24C36_GB40 = R24C36_GBO1;
assign R24C37_GB40 = R24C36_GBO1;
assign R24C38_GB40 = R24C36_GBO1;
assign R25C35_GB40 = R25C36_GBO1;
assign R25C36_GB40 = R25C36_GBO1;
assign R25C37_GB40 = R25C36_GBO1;
assign R25C38_GB40 = R25C36_GBO1;
assign R26C35_GB40 = R26C36_GBO1;
assign R26C36_GB40 = R26C36_GBO1;
assign R26C37_GB40 = R26C36_GBO1;
assign R26C38_GB40 = R26C36_GBO1;
assign R27C35_GB40 = R27C36_GBO1;
assign R27C36_GB40 = R27C36_GBO1;
assign R27C37_GB40 = R27C36_GBO1;
assign R27C38_GB40 = R27C36_GBO1;
assign R11C41_GB40 = R11C40_GBO1;
assign R11C42_GB40 = R11C40_GBO1;
assign R11C39_GB40 = R11C40_GBO1;
assign R11C40_GB40 = R11C40_GBO1;
assign R12C41_GB40 = R12C40_GBO1;
assign R12C42_GB40 = R12C40_GBO1;
assign R12C39_GB40 = R12C40_GBO1;
assign R12C40_GB40 = R12C40_GBO1;
assign R13C41_GB40 = R13C40_GBO1;
assign R13C42_GB40 = R13C40_GBO1;
assign R13C39_GB40 = R13C40_GBO1;
assign R13C40_GB40 = R13C40_GBO1;
assign R14C41_GB40 = R14C40_GBO1;
assign R14C42_GB40 = R14C40_GBO1;
assign R14C39_GB40 = R14C40_GBO1;
assign R14C40_GB40 = R14C40_GBO1;
assign R15C41_GB40 = R15C40_GBO1;
assign R15C42_GB40 = R15C40_GBO1;
assign R15C39_GB40 = R15C40_GBO1;
assign R15C40_GB40 = R15C40_GBO1;
assign R16C41_GB40 = R16C40_GBO1;
assign R16C42_GB40 = R16C40_GBO1;
assign R16C39_GB40 = R16C40_GBO1;
assign R16C40_GB40 = R16C40_GBO1;
assign R17C41_GB40 = R17C40_GBO1;
assign R17C42_GB40 = R17C40_GBO1;
assign R17C39_GB40 = R17C40_GBO1;
assign R17C40_GB40 = R17C40_GBO1;
assign R18C41_GB40 = R18C40_GBO1;
assign R18C42_GB40 = R18C40_GBO1;
assign R18C39_GB40 = R18C40_GBO1;
assign R18C40_GB40 = R18C40_GBO1;
assign R20C41_GB40 = R20C40_GBO1;
assign R20C42_GB40 = R20C40_GBO1;
assign R20C39_GB40 = R20C40_GBO1;
assign R20C40_GB40 = R20C40_GBO1;
assign R21C41_GB40 = R21C40_GBO1;
assign R21C42_GB40 = R21C40_GBO1;
assign R21C39_GB40 = R21C40_GBO1;
assign R21C40_GB40 = R21C40_GBO1;
assign R22C41_GB40 = R22C40_GBO1;
assign R22C42_GB40 = R22C40_GBO1;
assign R22C39_GB40 = R22C40_GBO1;
assign R22C40_GB40 = R22C40_GBO1;
assign R23C41_GB40 = R23C40_GBO1;
assign R23C42_GB40 = R23C40_GBO1;
assign R23C39_GB40 = R23C40_GBO1;
assign R23C40_GB40 = R23C40_GBO1;
assign R24C41_GB40 = R24C40_GBO1;
assign R24C42_GB40 = R24C40_GBO1;
assign R24C39_GB40 = R24C40_GBO1;
assign R24C40_GB40 = R24C40_GBO1;
assign R25C41_GB40 = R25C40_GBO1;
assign R25C42_GB40 = R25C40_GBO1;
assign R25C39_GB40 = R25C40_GBO1;
assign R25C40_GB40 = R25C40_GBO1;
assign R26C41_GB40 = R26C40_GBO1;
assign R26C42_GB40 = R26C40_GBO1;
assign R26C39_GB40 = R26C40_GBO1;
assign R26C40_GB40 = R26C40_GBO1;
assign R27C41_GB40 = R27C40_GBO1;
assign R27C42_GB40 = R27C40_GBO1;
assign R27C39_GB40 = R27C40_GBO1;
assign R27C40_GB40 = R27C40_GBO1;
assign R11C43_GB40 = R11C44_GBO1;
assign R11C44_GB40 = R11C44_GBO1;
assign R11C45_GB40 = R11C44_GBO1;
assign R11C46_GB40 = R11C44_GBO1;
assign R12C43_GB40 = R12C44_GBO1;
assign R12C44_GB40 = R12C44_GBO1;
assign R12C45_GB40 = R12C44_GBO1;
assign R12C46_GB40 = R12C44_GBO1;
assign R13C43_GB40 = R13C44_GBO1;
assign R13C44_GB40 = R13C44_GBO1;
assign R13C45_GB40 = R13C44_GBO1;
assign R13C46_GB40 = R13C44_GBO1;
assign R14C43_GB40 = R14C44_GBO1;
assign R14C44_GB40 = R14C44_GBO1;
assign R14C45_GB40 = R14C44_GBO1;
assign R14C46_GB40 = R14C44_GBO1;
assign R15C43_GB40 = R15C44_GBO1;
assign R15C44_GB40 = R15C44_GBO1;
assign R15C45_GB40 = R15C44_GBO1;
assign R15C46_GB40 = R15C44_GBO1;
assign R16C43_GB40 = R16C44_GBO1;
assign R16C44_GB40 = R16C44_GBO1;
assign R16C45_GB40 = R16C44_GBO1;
assign R16C46_GB40 = R16C44_GBO1;
assign R17C43_GB40 = R17C44_GBO1;
assign R17C44_GB40 = R17C44_GBO1;
assign R17C45_GB40 = R17C44_GBO1;
assign R17C46_GB40 = R17C44_GBO1;
assign R18C43_GB40 = R18C44_GBO1;
assign R18C44_GB40 = R18C44_GBO1;
assign R18C45_GB40 = R18C44_GBO1;
assign R18C46_GB40 = R18C44_GBO1;
assign R20C43_GB40 = R20C44_GBO1;
assign R20C44_GB40 = R20C44_GBO1;
assign R20C45_GB40 = R20C44_GBO1;
assign R20C46_GB40 = R20C44_GBO1;
assign R21C43_GB40 = R21C44_GBO1;
assign R21C44_GB40 = R21C44_GBO1;
assign R21C45_GB40 = R21C44_GBO1;
assign R21C46_GB40 = R21C44_GBO1;
assign R22C43_GB40 = R22C44_GBO1;
assign R22C44_GB40 = R22C44_GBO1;
assign R22C45_GB40 = R22C44_GBO1;
assign R22C46_GB40 = R22C44_GBO1;
assign R23C43_GB40 = R23C44_GBO1;
assign R23C44_GB40 = R23C44_GBO1;
assign R23C45_GB40 = R23C44_GBO1;
assign R23C46_GB40 = R23C44_GBO1;
assign R24C43_GB40 = R24C44_GBO1;
assign R24C44_GB40 = R24C44_GBO1;
assign R24C45_GB40 = R24C44_GBO1;
assign R24C46_GB40 = R24C44_GBO1;
assign R25C43_GB40 = R25C44_GBO1;
assign R25C44_GB40 = R25C44_GBO1;
assign R25C45_GB40 = R25C44_GBO1;
assign R25C46_GB40 = R25C44_GBO1;
assign R26C43_GB40 = R26C44_GBO1;
assign R26C44_GB40 = R26C44_GBO1;
assign R26C45_GB40 = R26C44_GBO1;
assign R26C46_GB40 = R26C44_GBO1;
assign R27C43_GB40 = R27C44_GBO1;
assign R27C44_GB40 = R27C44_GBO1;
assign R27C45_GB40 = R27C44_GBO1;
assign R27C46_GB40 = R27C44_GBO1;
assign R11C33_GB50 = R11C31_GBO1;
assign R11C29_GB50 = R11C31_GBO1;
assign R11C30_GB50 = R11C31_GBO1;
assign R11C31_GB50 = R11C31_GBO1;
assign R11C32_GB50 = R11C31_GBO1;
assign R12C33_GB50 = R12C31_GBO1;
assign R12C29_GB50 = R12C31_GBO1;
assign R12C30_GB50 = R12C31_GBO1;
assign R12C31_GB50 = R12C31_GBO1;
assign R12C32_GB50 = R12C31_GBO1;
assign R13C33_GB50 = R13C31_GBO1;
assign R13C29_GB50 = R13C31_GBO1;
assign R13C30_GB50 = R13C31_GBO1;
assign R13C31_GB50 = R13C31_GBO1;
assign R13C32_GB50 = R13C31_GBO1;
assign R14C33_GB50 = R14C31_GBO1;
assign R14C29_GB50 = R14C31_GBO1;
assign R14C30_GB50 = R14C31_GBO1;
assign R14C31_GB50 = R14C31_GBO1;
assign R14C32_GB50 = R14C31_GBO1;
assign R15C33_GB50 = R15C31_GBO1;
assign R15C29_GB50 = R15C31_GBO1;
assign R15C30_GB50 = R15C31_GBO1;
assign R15C31_GB50 = R15C31_GBO1;
assign R15C32_GB50 = R15C31_GBO1;
assign R16C33_GB50 = R16C31_GBO1;
assign R16C29_GB50 = R16C31_GBO1;
assign R16C30_GB50 = R16C31_GBO1;
assign R16C31_GB50 = R16C31_GBO1;
assign R16C32_GB50 = R16C31_GBO1;
assign R17C33_GB50 = R17C31_GBO1;
assign R17C29_GB50 = R17C31_GBO1;
assign R17C30_GB50 = R17C31_GBO1;
assign R17C31_GB50 = R17C31_GBO1;
assign R17C32_GB50 = R17C31_GBO1;
assign R18C33_GB50 = R18C31_GBO1;
assign R18C29_GB50 = R18C31_GBO1;
assign R18C30_GB50 = R18C31_GBO1;
assign R18C31_GB50 = R18C31_GBO1;
assign R18C32_GB50 = R18C31_GBO1;
assign R20C33_GB50 = R20C31_GBO1;
assign R20C29_GB50 = R20C31_GBO1;
assign R20C30_GB50 = R20C31_GBO1;
assign R20C31_GB50 = R20C31_GBO1;
assign R20C32_GB50 = R20C31_GBO1;
assign R21C33_GB50 = R21C31_GBO1;
assign R21C29_GB50 = R21C31_GBO1;
assign R21C30_GB50 = R21C31_GBO1;
assign R21C31_GB50 = R21C31_GBO1;
assign R21C32_GB50 = R21C31_GBO1;
assign R22C33_GB50 = R22C31_GBO1;
assign R22C29_GB50 = R22C31_GBO1;
assign R22C30_GB50 = R22C31_GBO1;
assign R22C31_GB50 = R22C31_GBO1;
assign R22C32_GB50 = R22C31_GBO1;
assign R23C33_GB50 = R23C31_GBO1;
assign R23C29_GB50 = R23C31_GBO1;
assign R23C30_GB50 = R23C31_GBO1;
assign R23C31_GB50 = R23C31_GBO1;
assign R23C32_GB50 = R23C31_GBO1;
assign R24C33_GB50 = R24C31_GBO1;
assign R24C29_GB50 = R24C31_GBO1;
assign R24C30_GB50 = R24C31_GBO1;
assign R24C31_GB50 = R24C31_GBO1;
assign R24C32_GB50 = R24C31_GBO1;
assign R25C33_GB50 = R25C31_GBO1;
assign R25C29_GB50 = R25C31_GBO1;
assign R25C30_GB50 = R25C31_GBO1;
assign R25C31_GB50 = R25C31_GBO1;
assign R25C32_GB50 = R25C31_GBO1;
assign R26C33_GB50 = R26C31_GBO1;
assign R26C29_GB50 = R26C31_GBO1;
assign R26C30_GB50 = R26C31_GBO1;
assign R26C31_GB50 = R26C31_GBO1;
assign R26C32_GB50 = R26C31_GBO1;
assign R27C33_GB50 = R27C31_GBO1;
assign R27C29_GB50 = R27C31_GBO1;
assign R27C30_GB50 = R27C31_GBO1;
assign R27C31_GB50 = R27C31_GBO1;
assign R27C32_GB50 = R27C31_GBO1;
assign R11C34_GB50 = R11C35_GBO1;
assign R11C35_GB50 = R11C35_GBO1;
assign R11C36_GB50 = R11C35_GBO1;
assign R11C37_GB50 = R11C35_GBO1;
assign R12C34_GB50 = R12C35_GBO1;
assign R12C35_GB50 = R12C35_GBO1;
assign R12C36_GB50 = R12C35_GBO1;
assign R12C37_GB50 = R12C35_GBO1;
assign R13C34_GB50 = R13C35_GBO1;
assign R13C35_GB50 = R13C35_GBO1;
assign R13C36_GB50 = R13C35_GBO1;
assign R13C37_GB50 = R13C35_GBO1;
assign R14C34_GB50 = R14C35_GBO1;
assign R14C35_GB50 = R14C35_GBO1;
assign R14C36_GB50 = R14C35_GBO1;
assign R14C37_GB50 = R14C35_GBO1;
assign R15C34_GB50 = R15C35_GBO1;
assign R15C35_GB50 = R15C35_GBO1;
assign R15C36_GB50 = R15C35_GBO1;
assign R15C37_GB50 = R15C35_GBO1;
assign R16C34_GB50 = R16C35_GBO1;
assign R16C35_GB50 = R16C35_GBO1;
assign R16C36_GB50 = R16C35_GBO1;
assign R16C37_GB50 = R16C35_GBO1;
assign R17C34_GB50 = R17C35_GBO1;
assign R17C35_GB50 = R17C35_GBO1;
assign R17C36_GB50 = R17C35_GBO1;
assign R17C37_GB50 = R17C35_GBO1;
assign R18C34_GB50 = R18C35_GBO1;
assign R18C35_GB50 = R18C35_GBO1;
assign R18C36_GB50 = R18C35_GBO1;
assign R18C37_GB50 = R18C35_GBO1;
assign R20C34_GB50 = R20C35_GBO1;
assign R20C35_GB50 = R20C35_GBO1;
assign R20C36_GB50 = R20C35_GBO1;
assign R20C37_GB50 = R20C35_GBO1;
assign R21C34_GB50 = R21C35_GBO1;
assign R21C35_GB50 = R21C35_GBO1;
assign R21C36_GB50 = R21C35_GBO1;
assign R21C37_GB50 = R21C35_GBO1;
assign R22C34_GB50 = R22C35_GBO1;
assign R22C35_GB50 = R22C35_GBO1;
assign R22C36_GB50 = R22C35_GBO1;
assign R22C37_GB50 = R22C35_GBO1;
assign R23C34_GB50 = R23C35_GBO1;
assign R23C35_GB50 = R23C35_GBO1;
assign R23C36_GB50 = R23C35_GBO1;
assign R23C37_GB50 = R23C35_GBO1;
assign R24C34_GB50 = R24C35_GBO1;
assign R24C35_GB50 = R24C35_GBO1;
assign R24C36_GB50 = R24C35_GBO1;
assign R24C37_GB50 = R24C35_GBO1;
assign R25C34_GB50 = R25C35_GBO1;
assign R25C35_GB50 = R25C35_GBO1;
assign R25C36_GB50 = R25C35_GBO1;
assign R25C37_GB50 = R25C35_GBO1;
assign R26C34_GB50 = R26C35_GBO1;
assign R26C35_GB50 = R26C35_GBO1;
assign R26C36_GB50 = R26C35_GBO1;
assign R26C37_GB50 = R26C35_GBO1;
assign R27C34_GB50 = R27C35_GBO1;
assign R27C35_GB50 = R27C35_GBO1;
assign R27C36_GB50 = R27C35_GBO1;
assign R27C37_GB50 = R27C35_GBO1;
assign R11C41_GB50 = R11C39_GBO1;
assign R11C38_GB50 = R11C39_GBO1;
assign R11C39_GB50 = R11C39_GBO1;
assign R11C40_GB50 = R11C39_GBO1;
assign R12C41_GB50 = R12C39_GBO1;
assign R12C38_GB50 = R12C39_GBO1;
assign R12C39_GB50 = R12C39_GBO1;
assign R12C40_GB50 = R12C39_GBO1;
assign R13C41_GB50 = R13C39_GBO1;
assign R13C38_GB50 = R13C39_GBO1;
assign R13C39_GB50 = R13C39_GBO1;
assign R13C40_GB50 = R13C39_GBO1;
assign R14C41_GB50 = R14C39_GBO1;
assign R14C38_GB50 = R14C39_GBO1;
assign R14C39_GB50 = R14C39_GBO1;
assign R14C40_GB50 = R14C39_GBO1;
assign R15C41_GB50 = R15C39_GBO1;
assign R15C38_GB50 = R15C39_GBO1;
assign R15C39_GB50 = R15C39_GBO1;
assign R15C40_GB50 = R15C39_GBO1;
assign R16C41_GB50 = R16C39_GBO1;
assign R16C38_GB50 = R16C39_GBO1;
assign R16C39_GB50 = R16C39_GBO1;
assign R16C40_GB50 = R16C39_GBO1;
assign R17C41_GB50 = R17C39_GBO1;
assign R17C38_GB50 = R17C39_GBO1;
assign R17C39_GB50 = R17C39_GBO1;
assign R17C40_GB50 = R17C39_GBO1;
assign R18C41_GB50 = R18C39_GBO1;
assign R18C38_GB50 = R18C39_GBO1;
assign R18C39_GB50 = R18C39_GBO1;
assign R18C40_GB50 = R18C39_GBO1;
assign R20C41_GB50 = R20C39_GBO1;
assign R20C38_GB50 = R20C39_GBO1;
assign R20C39_GB50 = R20C39_GBO1;
assign R20C40_GB50 = R20C39_GBO1;
assign R21C41_GB50 = R21C39_GBO1;
assign R21C38_GB50 = R21C39_GBO1;
assign R21C39_GB50 = R21C39_GBO1;
assign R21C40_GB50 = R21C39_GBO1;
assign R22C41_GB50 = R22C39_GBO1;
assign R22C38_GB50 = R22C39_GBO1;
assign R22C39_GB50 = R22C39_GBO1;
assign R22C40_GB50 = R22C39_GBO1;
assign R23C41_GB50 = R23C39_GBO1;
assign R23C38_GB50 = R23C39_GBO1;
assign R23C39_GB50 = R23C39_GBO1;
assign R23C40_GB50 = R23C39_GBO1;
assign R24C41_GB50 = R24C39_GBO1;
assign R24C38_GB50 = R24C39_GBO1;
assign R24C39_GB50 = R24C39_GBO1;
assign R24C40_GB50 = R24C39_GBO1;
assign R25C41_GB50 = R25C39_GBO1;
assign R25C38_GB50 = R25C39_GBO1;
assign R25C39_GB50 = R25C39_GBO1;
assign R25C40_GB50 = R25C39_GBO1;
assign R26C41_GB50 = R26C39_GBO1;
assign R26C38_GB50 = R26C39_GBO1;
assign R26C39_GB50 = R26C39_GBO1;
assign R26C40_GB50 = R26C39_GBO1;
assign R27C41_GB50 = R27C39_GBO1;
assign R27C38_GB50 = R27C39_GBO1;
assign R27C39_GB50 = R27C39_GBO1;
assign R27C40_GB50 = R27C39_GBO1;
assign R11C42_GB50 = R11C43_GBO1;
assign R11C43_GB50 = R11C43_GBO1;
assign R11C44_GB50 = R11C43_GBO1;
assign R11C45_GB50 = R11C43_GBO1;
assign R11C46_GB50 = R11C43_GBO1;
assign R12C42_GB50 = R12C43_GBO1;
assign R12C43_GB50 = R12C43_GBO1;
assign R12C44_GB50 = R12C43_GBO1;
assign R12C45_GB50 = R12C43_GBO1;
assign R12C46_GB50 = R12C43_GBO1;
assign R13C42_GB50 = R13C43_GBO1;
assign R13C43_GB50 = R13C43_GBO1;
assign R13C44_GB50 = R13C43_GBO1;
assign R13C45_GB50 = R13C43_GBO1;
assign R13C46_GB50 = R13C43_GBO1;
assign R14C42_GB50 = R14C43_GBO1;
assign R14C43_GB50 = R14C43_GBO1;
assign R14C44_GB50 = R14C43_GBO1;
assign R14C45_GB50 = R14C43_GBO1;
assign R14C46_GB50 = R14C43_GBO1;
assign R15C42_GB50 = R15C43_GBO1;
assign R15C43_GB50 = R15C43_GBO1;
assign R15C44_GB50 = R15C43_GBO1;
assign R15C45_GB50 = R15C43_GBO1;
assign R15C46_GB50 = R15C43_GBO1;
assign R16C42_GB50 = R16C43_GBO1;
assign R16C43_GB50 = R16C43_GBO1;
assign R16C44_GB50 = R16C43_GBO1;
assign R16C45_GB50 = R16C43_GBO1;
assign R16C46_GB50 = R16C43_GBO1;
assign R17C42_GB50 = R17C43_GBO1;
assign R17C43_GB50 = R17C43_GBO1;
assign R17C44_GB50 = R17C43_GBO1;
assign R17C45_GB50 = R17C43_GBO1;
assign R17C46_GB50 = R17C43_GBO1;
assign R18C42_GB50 = R18C43_GBO1;
assign R18C43_GB50 = R18C43_GBO1;
assign R18C44_GB50 = R18C43_GBO1;
assign R18C45_GB50 = R18C43_GBO1;
assign R18C46_GB50 = R18C43_GBO1;
assign R20C42_GB50 = R20C43_GBO1;
assign R20C43_GB50 = R20C43_GBO1;
assign R20C44_GB50 = R20C43_GBO1;
assign R20C45_GB50 = R20C43_GBO1;
assign R20C46_GB50 = R20C43_GBO1;
assign R21C42_GB50 = R21C43_GBO1;
assign R21C43_GB50 = R21C43_GBO1;
assign R21C44_GB50 = R21C43_GBO1;
assign R21C45_GB50 = R21C43_GBO1;
assign R21C46_GB50 = R21C43_GBO1;
assign R22C42_GB50 = R22C43_GBO1;
assign R22C43_GB50 = R22C43_GBO1;
assign R22C44_GB50 = R22C43_GBO1;
assign R22C45_GB50 = R22C43_GBO1;
assign R22C46_GB50 = R22C43_GBO1;
assign R23C42_GB50 = R23C43_GBO1;
assign R23C43_GB50 = R23C43_GBO1;
assign R23C44_GB50 = R23C43_GBO1;
assign R23C45_GB50 = R23C43_GBO1;
assign R23C46_GB50 = R23C43_GBO1;
assign R24C42_GB50 = R24C43_GBO1;
assign R24C43_GB50 = R24C43_GBO1;
assign R24C44_GB50 = R24C43_GBO1;
assign R24C45_GB50 = R24C43_GBO1;
assign R24C46_GB50 = R24C43_GBO1;
assign R25C42_GB50 = R25C43_GBO1;
assign R25C43_GB50 = R25C43_GBO1;
assign R25C44_GB50 = R25C43_GBO1;
assign R25C45_GB50 = R25C43_GBO1;
assign R25C46_GB50 = R25C43_GBO1;
assign R26C42_GB50 = R26C43_GBO1;
assign R26C43_GB50 = R26C43_GBO1;
assign R26C44_GB50 = R26C43_GBO1;
assign R26C45_GB50 = R26C43_GBO1;
assign R26C46_GB50 = R26C43_GBO1;
assign R27C42_GB50 = R27C43_GBO1;
assign R27C43_GB50 = R27C43_GBO1;
assign R27C44_GB50 = R27C43_GBO1;
assign R27C45_GB50 = R27C43_GBO1;
assign R27C46_GB50 = R27C43_GBO1;
assign R11C29_GB60 = R11C30_GBO1;
assign R11C30_GB60 = R11C30_GBO1;
assign R11C31_GB60 = R11C30_GBO1;
assign R11C32_GB60 = R11C30_GBO1;
assign R12C29_GB60 = R12C30_GBO1;
assign R12C30_GB60 = R12C30_GBO1;
assign R12C31_GB60 = R12C30_GBO1;
assign R12C32_GB60 = R12C30_GBO1;
assign R13C29_GB60 = R13C30_GBO1;
assign R13C30_GB60 = R13C30_GBO1;
assign R13C31_GB60 = R13C30_GBO1;
assign R13C32_GB60 = R13C30_GBO1;
assign R14C29_GB60 = R14C30_GBO1;
assign R14C30_GB60 = R14C30_GBO1;
assign R14C31_GB60 = R14C30_GBO1;
assign R14C32_GB60 = R14C30_GBO1;
assign R15C29_GB60 = R15C30_GBO1;
assign R15C30_GB60 = R15C30_GBO1;
assign R15C31_GB60 = R15C30_GBO1;
assign R15C32_GB60 = R15C30_GBO1;
assign R16C29_GB60 = R16C30_GBO1;
assign R16C30_GB60 = R16C30_GBO1;
assign R16C31_GB60 = R16C30_GBO1;
assign R16C32_GB60 = R16C30_GBO1;
assign R17C29_GB60 = R17C30_GBO1;
assign R17C30_GB60 = R17C30_GBO1;
assign R17C31_GB60 = R17C30_GBO1;
assign R17C32_GB60 = R17C30_GBO1;
assign R18C29_GB60 = R18C30_GBO1;
assign R18C30_GB60 = R18C30_GBO1;
assign R18C31_GB60 = R18C30_GBO1;
assign R18C32_GB60 = R18C30_GBO1;
assign R20C29_GB60 = R20C30_GBO1;
assign R20C30_GB60 = R20C30_GBO1;
assign R20C31_GB60 = R20C30_GBO1;
assign R20C32_GB60 = R20C30_GBO1;
assign R21C29_GB60 = R21C30_GBO1;
assign R21C30_GB60 = R21C30_GBO1;
assign R21C31_GB60 = R21C30_GBO1;
assign R21C32_GB60 = R21C30_GBO1;
assign R22C29_GB60 = R22C30_GBO1;
assign R22C30_GB60 = R22C30_GBO1;
assign R22C31_GB60 = R22C30_GBO1;
assign R22C32_GB60 = R22C30_GBO1;
assign R23C29_GB60 = R23C30_GBO1;
assign R23C30_GB60 = R23C30_GBO1;
assign R23C31_GB60 = R23C30_GBO1;
assign R23C32_GB60 = R23C30_GBO1;
assign R24C29_GB60 = R24C30_GBO1;
assign R24C30_GB60 = R24C30_GBO1;
assign R24C31_GB60 = R24C30_GBO1;
assign R24C32_GB60 = R24C30_GBO1;
assign R25C29_GB60 = R25C30_GBO1;
assign R25C30_GB60 = R25C30_GBO1;
assign R25C31_GB60 = R25C30_GBO1;
assign R25C32_GB60 = R25C30_GBO1;
assign R26C29_GB60 = R26C30_GBO1;
assign R26C30_GB60 = R26C30_GBO1;
assign R26C31_GB60 = R26C30_GBO1;
assign R26C32_GB60 = R26C30_GBO1;
assign R27C29_GB60 = R27C30_GBO1;
assign R27C30_GB60 = R27C30_GBO1;
assign R27C31_GB60 = R27C30_GBO1;
assign R27C32_GB60 = R27C30_GBO1;
assign R11C33_GB60 = R11C34_GBO1;
assign R11C34_GB60 = R11C34_GBO1;
assign R11C35_GB60 = R11C34_GBO1;
assign R11C36_GB60 = R11C34_GBO1;
assign R12C33_GB60 = R12C34_GBO1;
assign R12C34_GB60 = R12C34_GBO1;
assign R12C35_GB60 = R12C34_GBO1;
assign R12C36_GB60 = R12C34_GBO1;
assign R13C33_GB60 = R13C34_GBO1;
assign R13C34_GB60 = R13C34_GBO1;
assign R13C35_GB60 = R13C34_GBO1;
assign R13C36_GB60 = R13C34_GBO1;
assign R14C33_GB60 = R14C34_GBO1;
assign R14C34_GB60 = R14C34_GBO1;
assign R14C35_GB60 = R14C34_GBO1;
assign R14C36_GB60 = R14C34_GBO1;
assign R15C33_GB60 = R15C34_GBO1;
assign R15C34_GB60 = R15C34_GBO1;
assign R15C35_GB60 = R15C34_GBO1;
assign R15C36_GB60 = R15C34_GBO1;
assign R16C33_GB60 = R16C34_GBO1;
assign R16C34_GB60 = R16C34_GBO1;
assign R16C35_GB60 = R16C34_GBO1;
assign R16C36_GB60 = R16C34_GBO1;
assign R17C33_GB60 = R17C34_GBO1;
assign R17C34_GB60 = R17C34_GBO1;
assign R17C35_GB60 = R17C34_GBO1;
assign R17C36_GB60 = R17C34_GBO1;
assign R18C33_GB60 = R18C34_GBO1;
assign R18C34_GB60 = R18C34_GBO1;
assign R18C35_GB60 = R18C34_GBO1;
assign R18C36_GB60 = R18C34_GBO1;
assign R20C33_GB60 = R20C34_GBO1;
assign R20C34_GB60 = R20C34_GBO1;
assign R20C35_GB60 = R20C34_GBO1;
assign R20C36_GB60 = R20C34_GBO1;
assign R21C33_GB60 = R21C34_GBO1;
assign R21C34_GB60 = R21C34_GBO1;
assign R21C35_GB60 = R21C34_GBO1;
assign R21C36_GB60 = R21C34_GBO1;
assign R22C33_GB60 = R22C34_GBO1;
assign R22C34_GB60 = R22C34_GBO1;
assign R22C35_GB60 = R22C34_GBO1;
assign R22C36_GB60 = R22C34_GBO1;
assign R23C33_GB60 = R23C34_GBO1;
assign R23C34_GB60 = R23C34_GBO1;
assign R23C35_GB60 = R23C34_GBO1;
assign R23C36_GB60 = R23C34_GBO1;
assign R24C33_GB60 = R24C34_GBO1;
assign R24C34_GB60 = R24C34_GBO1;
assign R24C35_GB60 = R24C34_GBO1;
assign R24C36_GB60 = R24C34_GBO1;
assign R25C33_GB60 = R25C34_GBO1;
assign R25C34_GB60 = R25C34_GBO1;
assign R25C35_GB60 = R25C34_GBO1;
assign R25C36_GB60 = R25C34_GBO1;
assign R26C33_GB60 = R26C34_GBO1;
assign R26C34_GB60 = R26C34_GBO1;
assign R26C35_GB60 = R26C34_GBO1;
assign R26C36_GB60 = R26C34_GBO1;
assign R27C33_GB60 = R27C34_GBO1;
assign R27C34_GB60 = R27C34_GBO1;
assign R27C35_GB60 = R27C34_GBO1;
assign R27C36_GB60 = R27C34_GBO1;
assign R11C37_GB60 = R11C38_GBO1;
assign R11C38_GB60 = R11C38_GBO1;
assign R11C39_GB60 = R11C38_GBO1;
assign R11C40_GB60 = R11C38_GBO1;
assign R12C37_GB60 = R12C38_GBO1;
assign R12C38_GB60 = R12C38_GBO1;
assign R12C39_GB60 = R12C38_GBO1;
assign R12C40_GB60 = R12C38_GBO1;
assign R13C37_GB60 = R13C38_GBO1;
assign R13C38_GB60 = R13C38_GBO1;
assign R13C39_GB60 = R13C38_GBO1;
assign R13C40_GB60 = R13C38_GBO1;
assign R14C37_GB60 = R14C38_GBO1;
assign R14C38_GB60 = R14C38_GBO1;
assign R14C39_GB60 = R14C38_GBO1;
assign R14C40_GB60 = R14C38_GBO1;
assign R15C37_GB60 = R15C38_GBO1;
assign R15C38_GB60 = R15C38_GBO1;
assign R15C39_GB60 = R15C38_GBO1;
assign R15C40_GB60 = R15C38_GBO1;
assign R16C37_GB60 = R16C38_GBO1;
assign R16C38_GB60 = R16C38_GBO1;
assign R16C39_GB60 = R16C38_GBO1;
assign R16C40_GB60 = R16C38_GBO1;
assign R17C37_GB60 = R17C38_GBO1;
assign R17C38_GB60 = R17C38_GBO1;
assign R17C39_GB60 = R17C38_GBO1;
assign R17C40_GB60 = R17C38_GBO1;
assign R18C37_GB60 = R18C38_GBO1;
assign R18C38_GB60 = R18C38_GBO1;
assign R18C39_GB60 = R18C38_GBO1;
assign R18C40_GB60 = R18C38_GBO1;
assign R20C37_GB60 = R20C38_GBO1;
assign R20C38_GB60 = R20C38_GBO1;
assign R20C39_GB60 = R20C38_GBO1;
assign R20C40_GB60 = R20C38_GBO1;
assign R21C37_GB60 = R21C38_GBO1;
assign R21C38_GB60 = R21C38_GBO1;
assign R21C39_GB60 = R21C38_GBO1;
assign R21C40_GB60 = R21C38_GBO1;
assign R22C37_GB60 = R22C38_GBO1;
assign R22C38_GB60 = R22C38_GBO1;
assign R22C39_GB60 = R22C38_GBO1;
assign R22C40_GB60 = R22C38_GBO1;
assign R23C37_GB60 = R23C38_GBO1;
assign R23C38_GB60 = R23C38_GBO1;
assign R23C39_GB60 = R23C38_GBO1;
assign R23C40_GB60 = R23C38_GBO1;
assign R24C37_GB60 = R24C38_GBO1;
assign R24C38_GB60 = R24C38_GBO1;
assign R24C39_GB60 = R24C38_GBO1;
assign R24C40_GB60 = R24C38_GBO1;
assign R25C37_GB60 = R25C38_GBO1;
assign R25C38_GB60 = R25C38_GBO1;
assign R25C39_GB60 = R25C38_GBO1;
assign R25C40_GB60 = R25C38_GBO1;
assign R26C37_GB60 = R26C38_GBO1;
assign R26C38_GB60 = R26C38_GBO1;
assign R26C39_GB60 = R26C38_GBO1;
assign R26C40_GB60 = R26C38_GBO1;
assign R27C37_GB60 = R27C38_GBO1;
assign R27C38_GB60 = R27C38_GBO1;
assign R27C39_GB60 = R27C38_GBO1;
assign R27C40_GB60 = R27C38_GBO1;
assign R11C41_GB60 = R11C42_GBO1;
assign R11C42_GB60 = R11C42_GBO1;
assign R11C43_GB60 = R11C42_GBO1;
assign R11C44_GB60 = R11C42_GBO1;
assign R12C41_GB60 = R12C42_GBO1;
assign R12C42_GB60 = R12C42_GBO1;
assign R12C43_GB60 = R12C42_GBO1;
assign R12C44_GB60 = R12C42_GBO1;
assign R13C41_GB60 = R13C42_GBO1;
assign R13C42_GB60 = R13C42_GBO1;
assign R13C43_GB60 = R13C42_GBO1;
assign R13C44_GB60 = R13C42_GBO1;
assign R14C41_GB60 = R14C42_GBO1;
assign R14C42_GB60 = R14C42_GBO1;
assign R14C43_GB60 = R14C42_GBO1;
assign R14C44_GB60 = R14C42_GBO1;
assign R15C41_GB60 = R15C42_GBO1;
assign R15C42_GB60 = R15C42_GBO1;
assign R15C43_GB60 = R15C42_GBO1;
assign R15C44_GB60 = R15C42_GBO1;
assign R16C41_GB60 = R16C42_GBO1;
assign R16C42_GB60 = R16C42_GBO1;
assign R16C43_GB60 = R16C42_GBO1;
assign R16C44_GB60 = R16C42_GBO1;
assign R17C41_GB60 = R17C42_GBO1;
assign R17C42_GB60 = R17C42_GBO1;
assign R17C43_GB60 = R17C42_GBO1;
assign R17C44_GB60 = R17C42_GBO1;
assign R18C41_GB60 = R18C42_GBO1;
assign R18C42_GB60 = R18C42_GBO1;
assign R18C43_GB60 = R18C42_GBO1;
assign R18C44_GB60 = R18C42_GBO1;
assign R20C41_GB60 = R20C42_GBO1;
assign R20C42_GB60 = R20C42_GBO1;
assign R20C43_GB60 = R20C42_GBO1;
assign R20C44_GB60 = R20C42_GBO1;
assign R21C41_GB60 = R21C42_GBO1;
assign R21C42_GB60 = R21C42_GBO1;
assign R21C43_GB60 = R21C42_GBO1;
assign R21C44_GB60 = R21C42_GBO1;
assign R22C41_GB60 = R22C42_GBO1;
assign R22C42_GB60 = R22C42_GBO1;
assign R22C43_GB60 = R22C42_GBO1;
assign R22C44_GB60 = R22C42_GBO1;
assign R23C41_GB60 = R23C42_GBO1;
assign R23C42_GB60 = R23C42_GBO1;
assign R23C43_GB60 = R23C42_GBO1;
assign R23C44_GB60 = R23C42_GBO1;
assign R24C41_GB60 = R24C42_GBO1;
assign R24C42_GB60 = R24C42_GBO1;
assign R24C43_GB60 = R24C42_GBO1;
assign R24C44_GB60 = R24C42_GBO1;
assign R25C41_GB60 = R25C42_GBO1;
assign R25C42_GB60 = R25C42_GBO1;
assign R25C43_GB60 = R25C42_GBO1;
assign R25C44_GB60 = R25C42_GBO1;
assign R26C41_GB60 = R26C42_GBO1;
assign R26C42_GB60 = R26C42_GBO1;
assign R26C43_GB60 = R26C42_GBO1;
assign R26C44_GB60 = R26C42_GBO1;
assign R27C41_GB60 = R27C42_GBO1;
assign R27C42_GB60 = R27C42_GBO1;
assign R27C43_GB60 = R27C42_GBO1;
assign R27C44_GB60 = R27C42_GBO1;
assign R11C45_GB60 = R11C46_GBO1;
assign R11C46_GB60 = R11C46_GBO1;
assign R12C45_GB60 = R12C46_GBO1;
assign R12C46_GB60 = R12C46_GBO1;
assign R13C45_GB60 = R13C46_GBO1;
assign R13C46_GB60 = R13C46_GBO1;
assign R14C45_GB60 = R14C46_GBO1;
assign R14C46_GB60 = R14C46_GBO1;
assign R15C45_GB60 = R15C46_GBO1;
assign R15C46_GB60 = R15C46_GBO1;
assign R16C45_GB60 = R16C46_GBO1;
assign R16C46_GB60 = R16C46_GBO1;
assign R17C45_GB60 = R17C46_GBO1;
assign R17C46_GB60 = R17C46_GBO1;
assign R18C45_GB60 = R18C46_GBO1;
assign R18C46_GB60 = R18C46_GBO1;
assign R20C45_GB60 = R20C46_GBO1;
assign R20C46_GB60 = R20C46_GBO1;
assign R21C45_GB60 = R21C46_GBO1;
assign R21C46_GB60 = R21C46_GBO1;
assign R22C45_GB60 = R22C46_GBO1;
assign R22C46_GB60 = R22C46_GBO1;
assign R23C45_GB60 = R23C46_GBO1;
assign R23C46_GB60 = R23C46_GBO1;
assign R24C45_GB60 = R24C46_GBO1;
assign R24C46_GB60 = R24C46_GBO1;
assign R25C45_GB60 = R25C46_GBO1;
assign R25C46_GB60 = R25C46_GBO1;
assign R26C45_GB60 = R26C46_GBO1;
assign R26C46_GB60 = R26C46_GBO1;
assign R27C45_GB60 = R27C46_GBO1;
assign R27C46_GB60 = R27C46_GBO1;
assign R11C29_GB70 = R11C29_GBO1;
assign R11C30_GB70 = R11C29_GBO1;
assign R11C31_GB70 = R11C29_GBO1;
assign R12C29_GB70 = R12C29_GBO1;
assign R12C30_GB70 = R12C29_GBO1;
assign R12C31_GB70 = R12C29_GBO1;
assign R13C29_GB70 = R13C29_GBO1;
assign R13C30_GB70 = R13C29_GBO1;
assign R13C31_GB70 = R13C29_GBO1;
assign R14C29_GB70 = R14C29_GBO1;
assign R14C30_GB70 = R14C29_GBO1;
assign R14C31_GB70 = R14C29_GBO1;
assign R15C29_GB70 = R15C29_GBO1;
assign R15C30_GB70 = R15C29_GBO1;
assign R15C31_GB70 = R15C29_GBO1;
assign R16C29_GB70 = R16C29_GBO1;
assign R16C30_GB70 = R16C29_GBO1;
assign R16C31_GB70 = R16C29_GBO1;
assign R17C29_GB70 = R17C29_GBO1;
assign R17C30_GB70 = R17C29_GBO1;
assign R17C31_GB70 = R17C29_GBO1;
assign R18C29_GB70 = R18C29_GBO1;
assign R18C30_GB70 = R18C29_GBO1;
assign R18C31_GB70 = R18C29_GBO1;
assign R20C29_GB70 = R20C29_GBO1;
assign R20C30_GB70 = R20C29_GBO1;
assign R20C31_GB70 = R20C29_GBO1;
assign R21C29_GB70 = R21C29_GBO1;
assign R21C30_GB70 = R21C29_GBO1;
assign R21C31_GB70 = R21C29_GBO1;
assign R22C29_GB70 = R22C29_GBO1;
assign R22C30_GB70 = R22C29_GBO1;
assign R22C31_GB70 = R22C29_GBO1;
assign R23C29_GB70 = R23C29_GBO1;
assign R23C30_GB70 = R23C29_GBO1;
assign R23C31_GB70 = R23C29_GBO1;
assign R24C29_GB70 = R24C29_GBO1;
assign R24C30_GB70 = R24C29_GBO1;
assign R24C31_GB70 = R24C29_GBO1;
assign R25C29_GB70 = R25C29_GBO1;
assign R25C30_GB70 = R25C29_GBO1;
assign R25C31_GB70 = R25C29_GBO1;
assign R26C29_GB70 = R26C29_GBO1;
assign R26C30_GB70 = R26C29_GBO1;
assign R26C31_GB70 = R26C29_GBO1;
assign R27C29_GB70 = R27C29_GBO1;
assign R27C30_GB70 = R27C29_GBO1;
assign R27C31_GB70 = R27C29_GBO1;
assign R11C33_GB70 = R11C33_GBO1;
assign R11C34_GB70 = R11C33_GBO1;
assign R11C35_GB70 = R11C33_GBO1;
assign R11C32_GB70 = R11C33_GBO1;
assign R12C33_GB70 = R12C33_GBO1;
assign R12C34_GB70 = R12C33_GBO1;
assign R12C35_GB70 = R12C33_GBO1;
assign R12C32_GB70 = R12C33_GBO1;
assign R13C33_GB70 = R13C33_GBO1;
assign R13C34_GB70 = R13C33_GBO1;
assign R13C35_GB70 = R13C33_GBO1;
assign R13C32_GB70 = R13C33_GBO1;
assign R14C33_GB70 = R14C33_GBO1;
assign R14C34_GB70 = R14C33_GBO1;
assign R14C35_GB70 = R14C33_GBO1;
assign R14C32_GB70 = R14C33_GBO1;
assign R15C33_GB70 = R15C33_GBO1;
assign R15C34_GB70 = R15C33_GBO1;
assign R15C35_GB70 = R15C33_GBO1;
assign R15C32_GB70 = R15C33_GBO1;
assign R16C33_GB70 = R16C33_GBO1;
assign R16C34_GB70 = R16C33_GBO1;
assign R16C35_GB70 = R16C33_GBO1;
assign R16C32_GB70 = R16C33_GBO1;
assign R17C33_GB70 = R17C33_GBO1;
assign R17C34_GB70 = R17C33_GBO1;
assign R17C35_GB70 = R17C33_GBO1;
assign R17C32_GB70 = R17C33_GBO1;
assign R18C33_GB70 = R18C33_GBO1;
assign R18C34_GB70 = R18C33_GBO1;
assign R18C35_GB70 = R18C33_GBO1;
assign R18C32_GB70 = R18C33_GBO1;
assign R20C33_GB70 = R20C33_GBO1;
assign R20C34_GB70 = R20C33_GBO1;
assign R20C35_GB70 = R20C33_GBO1;
assign R20C32_GB70 = R20C33_GBO1;
assign R21C33_GB70 = R21C33_GBO1;
assign R21C34_GB70 = R21C33_GBO1;
assign R21C35_GB70 = R21C33_GBO1;
assign R21C32_GB70 = R21C33_GBO1;
assign R22C33_GB70 = R22C33_GBO1;
assign R22C34_GB70 = R22C33_GBO1;
assign R22C35_GB70 = R22C33_GBO1;
assign R22C32_GB70 = R22C33_GBO1;
assign R23C33_GB70 = R23C33_GBO1;
assign R23C34_GB70 = R23C33_GBO1;
assign R23C35_GB70 = R23C33_GBO1;
assign R23C32_GB70 = R23C33_GBO1;
assign R24C33_GB70 = R24C33_GBO1;
assign R24C34_GB70 = R24C33_GBO1;
assign R24C35_GB70 = R24C33_GBO1;
assign R24C32_GB70 = R24C33_GBO1;
assign R25C33_GB70 = R25C33_GBO1;
assign R25C34_GB70 = R25C33_GBO1;
assign R25C35_GB70 = R25C33_GBO1;
assign R25C32_GB70 = R25C33_GBO1;
assign R26C33_GB70 = R26C33_GBO1;
assign R26C34_GB70 = R26C33_GBO1;
assign R26C35_GB70 = R26C33_GBO1;
assign R26C32_GB70 = R26C33_GBO1;
assign R27C33_GB70 = R27C33_GBO1;
assign R27C34_GB70 = R27C33_GBO1;
assign R27C35_GB70 = R27C33_GBO1;
assign R27C32_GB70 = R27C33_GBO1;
assign R11C36_GB70 = R11C37_GBO1;
assign R11C37_GB70 = R11C37_GBO1;
assign R11C38_GB70 = R11C37_GBO1;
assign R11C39_GB70 = R11C37_GBO1;
assign R12C36_GB70 = R12C37_GBO1;
assign R12C37_GB70 = R12C37_GBO1;
assign R12C38_GB70 = R12C37_GBO1;
assign R12C39_GB70 = R12C37_GBO1;
assign R13C36_GB70 = R13C37_GBO1;
assign R13C37_GB70 = R13C37_GBO1;
assign R13C38_GB70 = R13C37_GBO1;
assign R13C39_GB70 = R13C37_GBO1;
assign R14C36_GB70 = R14C37_GBO1;
assign R14C37_GB70 = R14C37_GBO1;
assign R14C38_GB70 = R14C37_GBO1;
assign R14C39_GB70 = R14C37_GBO1;
assign R15C36_GB70 = R15C37_GBO1;
assign R15C37_GB70 = R15C37_GBO1;
assign R15C38_GB70 = R15C37_GBO1;
assign R15C39_GB70 = R15C37_GBO1;
assign R16C36_GB70 = R16C37_GBO1;
assign R16C37_GB70 = R16C37_GBO1;
assign R16C38_GB70 = R16C37_GBO1;
assign R16C39_GB70 = R16C37_GBO1;
assign R17C36_GB70 = R17C37_GBO1;
assign R17C37_GB70 = R17C37_GBO1;
assign R17C38_GB70 = R17C37_GBO1;
assign R17C39_GB70 = R17C37_GBO1;
assign R18C36_GB70 = R18C37_GBO1;
assign R18C37_GB70 = R18C37_GBO1;
assign R18C38_GB70 = R18C37_GBO1;
assign R18C39_GB70 = R18C37_GBO1;
assign R20C36_GB70 = R20C37_GBO1;
assign R20C37_GB70 = R20C37_GBO1;
assign R20C38_GB70 = R20C37_GBO1;
assign R20C39_GB70 = R20C37_GBO1;
assign R21C36_GB70 = R21C37_GBO1;
assign R21C37_GB70 = R21C37_GBO1;
assign R21C38_GB70 = R21C37_GBO1;
assign R21C39_GB70 = R21C37_GBO1;
assign R22C36_GB70 = R22C37_GBO1;
assign R22C37_GB70 = R22C37_GBO1;
assign R22C38_GB70 = R22C37_GBO1;
assign R22C39_GB70 = R22C37_GBO1;
assign R23C36_GB70 = R23C37_GBO1;
assign R23C37_GB70 = R23C37_GBO1;
assign R23C38_GB70 = R23C37_GBO1;
assign R23C39_GB70 = R23C37_GBO1;
assign R24C36_GB70 = R24C37_GBO1;
assign R24C37_GB70 = R24C37_GBO1;
assign R24C38_GB70 = R24C37_GBO1;
assign R24C39_GB70 = R24C37_GBO1;
assign R25C36_GB70 = R25C37_GBO1;
assign R25C37_GB70 = R25C37_GBO1;
assign R25C38_GB70 = R25C37_GBO1;
assign R25C39_GB70 = R25C37_GBO1;
assign R26C36_GB70 = R26C37_GBO1;
assign R26C37_GB70 = R26C37_GBO1;
assign R26C38_GB70 = R26C37_GBO1;
assign R26C39_GB70 = R26C37_GBO1;
assign R27C36_GB70 = R27C37_GBO1;
assign R27C37_GB70 = R27C37_GBO1;
assign R27C38_GB70 = R27C37_GBO1;
assign R27C39_GB70 = R27C37_GBO1;
assign R11C41_GB70 = R11C41_GBO1;
assign R11C42_GB70 = R11C41_GBO1;
assign R11C43_GB70 = R11C41_GBO1;
assign R11C40_GB70 = R11C41_GBO1;
assign R12C41_GB70 = R12C41_GBO1;
assign R12C42_GB70 = R12C41_GBO1;
assign R12C43_GB70 = R12C41_GBO1;
assign R12C40_GB70 = R12C41_GBO1;
assign R13C41_GB70 = R13C41_GBO1;
assign R13C42_GB70 = R13C41_GBO1;
assign R13C43_GB70 = R13C41_GBO1;
assign R13C40_GB70 = R13C41_GBO1;
assign R14C41_GB70 = R14C41_GBO1;
assign R14C42_GB70 = R14C41_GBO1;
assign R14C43_GB70 = R14C41_GBO1;
assign R14C40_GB70 = R14C41_GBO1;
assign R15C41_GB70 = R15C41_GBO1;
assign R15C42_GB70 = R15C41_GBO1;
assign R15C43_GB70 = R15C41_GBO1;
assign R15C40_GB70 = R15C41_GBO1;
assign R16C41_GB70 = R16C41_GBO1;
assign R16C42_GB70 = R16C41_GBO1;
assign R16C43_GB70 = R16C41_GBO1;
assign R16C40_GB70 = R16C41_GBO1;
assign R17C41_GB70 = R17C41_GBO1;
assign R17C42_GB70 = R17C41_GBO1;
assign R17C43_GB70 = R17C41_GBO1;
assign R17C40_GB70 = R17C41_GBO1;
assign R18C41_GB70 = R18C41_GBO1;
assign R18C42_GB70 = R18C41_GBO1;
assign R18C43_GB70 = R18C41_GBO1;
assign R18C40_GB70 = R18C41_GBO1;
assign R20C41_GB70 = R20C41_GBO1;
assign R20C42_GB70 = R20C41_GBO1;
assign R20C43_GB70 = R20C41_GBO1;
assign R20C40_GB70 = R20C41_GBO1;
assign R21C41_GB70 = R21C41_GBO1;
assign R21C42_GB70 = R21C41_GBO1;
assign R21C43_GB70 = R21C41_GBO1;
assign R21C40_GB70 = R21C41_GBO1;
assign R22C41_GB70 = R22C41_GBO1;
assign R22C42_GB70 = R22C41_GBO1;
assign R22C43_GB70 = R22C41_GBO1;
assign R22C40_GB70 = R22C41_GBO1;
assign R23C41_GB70 = R23C41_GBO1;
assign R23C42_GB70 = R23C41_GBO1;
assign R23C43_GB70 = R23C41_GBO1;
assign R23C40_GB70 = R23C41_GBO1;
assign R24C41_GB70 = R24C41_GBO1;
assign R24C42_GB70 = R24C41_GBO1;
assign R24C43_GB70 = R24C41_GBO1;
assign R24C40_GB70 = R24C41_GBO1;
assign R25C41_GB70 = R25C41_GBO1;
assign R25C42_GB70 = R25C41_GBO1;
assign R25C43_GB70 = R25C41_GBO1;
assign R25C40_GB70 = R25C41_GBO1;
assign R26C41_GB70 = R26C41_GBO1;
assign R26C42_GB70 = R26C41_GBO1;
assign R26C43_GB70 = R26C41_GBO1;
assign R26C40_GB70 = R26C41_GBO1;
assign R27C41_GB70 = R27C41_GBO1;
assign R27C42_GB70 = R27C41_GBO1;
assign R27C43_GB70 = R27C41_GBO1;
assign R27C40_GB70 = R27C41_GBO1;
assign R11C44_GB70 = R11C45_GBO1;
assign R11C45_GB70 = R11C45_GBO1;
assign R11C46_GB70 = R11C45_GBO1;
assign R12C44_GB70 = R12C45_GBO1;
assign R12C45_GB70 = R12C45_GBO1;
assign R12C46_GB70 = R12C45_GBO1;
assign R13C44_GB70 = R13C45_GBO1;
assign R13C45_GB70 = R13C45_GBO1;
assign R13C46_GB70 = R13C45_GBO1;
assign R14C44_GB70 = R14C45_GBO1;
assign R14C45_GB70 = R14C45_GBO1;
assign R14C46_GB70 = R14C45_GBO1;
assign R15C44_GB70 = R15C45_GBO1;
assign R15C45_GB70 = R15C45_GBO1;
assign R15C46_GB70 = R15C45_GBO1;
assign R16C44_GB70 = R16C45_GBO1;
assign R16C45_GB70 = R16C45_GBO1;
assign R16C46_GB70 = R16C45_GBO1;
assign R17C44_GB70 = R17C45_GBO1;
assign R17C45_GB70 = R17C45_GBO1;
assign R17C46_GB70 = R17C45_GBO1;
assign R18C44_GB70 = R18C45_GBO1;
assign R18C45_GB70 = R18C45_GBO1;
assign R18C46_GB70 = R18C45_GBO1;
assign R20C44_GB70 = R20C45_GBO1;
assign R20C45_GB70 = R20C45_GBO1;
assign R20C46_GB70 = R20C45_GBO1;
assign R21C44_GB70 = R21C45_GBO1;
assign R21C45_GB70 = R21C45_GBO1;
assign R21C46_GB70 = R21C45_GBO1;
assign R22C44_GB70 = R22C45_GBO1;
assign R22C45_GB70 = R22C45_GBO1;
assign R22C46_GB70 = R22C45_GBO1;
assign R23C44_GB70 = R23C45_GBO1;
assign R23C45_GB70 = R23C45_GBO1;
assign R23C46_GB70 = R23C45_GBO1;
assign R24C44_GB70 = R24C45_GBO1;
assign R24C45_GB70 = R24C45_GBO1;
assign R24C46_GB70 = R24C45_GBO1;
assign R25C44_GB70 = R25C45_GBO1;
assign R25C45_GB70 = R25C45_GBO1;
assign R25C46_GB70 = R25C45_GBO1;
assign R26C44_GB70 = R26C45_GBO1;
assign R26C45_GB70 = R26C45_GBO1;
assign R26C46_GB70 = R26C45_GBO1;
assign R27C44_GB70 = R27C45_GBO1;
assign R27C45_GB70 = R27C45_GBO1;
assign R27C46_GB70 = R27C45_GBO1;
assign R1C1_CLK0 = VCC;
assign R1C1_CLK1 = VCC;
assign R1C1_CLK2 = VCC;
assign R1C1_LSR0 = VCC;
assign R1C1_LSR1 = VCC;
assign R1C1_LSR2 = VCC;
assign R1C1_CE0 = VCC;
assign R1C1_CE1 = VCC;
assign R1C1_CE2 = VCC;
assign R1C1_SEL0 = VCC;
assign R1C1_SEL1 = VCC;
assign R1C1_SEL2 = VCC;
assign R1C1_SEL3 = VCC;
assign R1C1_SEL4 = VCC;
assign R1C1_SEL5 = VCC;
assign R1C1_SEL6 = VCC;
assign R1C1_SEL7 = VCC;
assign R1C1_C0 = R1C1_F4;
assign R1C1_C1 = R1C1_F4;
assign R1C1_C2 = R1C1_F4;
assign R1C1_C3 = R1C1_F4;
assign R1C1_A4 = R1C1_F7;
assign R1C1_A5 = R1C1_F7;
assign R1C1_A6 = R1C1_F5;
assign R1C1_A7 = R1C1_F5;
assign R1C1_N82 = R1C1_Q4;
assign R1C1_S82 = R1C1_Q4;
assign R1C1_E82 = R1C1_Q4;
assign R1C1_W82 = R1C1_Q4;
assign R1C1_A0 = R1C1_F5;
assign R1C1_A1 = R1C1_F5;
assign R1C1_A2 = R1C1_F5;
assign R1C1_A3 = R1C1_F5;
assign R1C1_C4 = R1C1_S22;
assign R1C1_C5 = R1C1_F6;
assign R1C1_C6 = R1C1_F4;
assign R1C1_C7 = R1C1_F4;
assign R1C1_N81 = R1C1_Q1;
assign R1C1_S81 = R1C1_Q1;
assign R1C1_E81 = R1C1_Q1;
assign R1C1_W81 = R1C1_Q1;
assign R1C1_N21 = R1C1_Q1;
assign R1C1_N22 = R1C1_Q2;
assign R1C1_S21 = R1C1_Q1;
assign R1C1_S22 = VCC;
assign R1C1_E21 = R1C1_Q1;
assign R1C1_E22 = R1C1_Q2;
assign R1C1_W21 = R1C1_Q1;
assign R1C1_W22 = R1C1_Q2;
assign R1C1_E80 = R1C1_Q0;
assign R1C1_W80 = R1C1_Q0;
assign R1C1_N25 = R1C1_Q5;
assign R1C1_N26 = R1C1_Q6;
assign R1C1_S25 = R1C1_Q5;
assign R1C1_S26 = R1C1_Q6;
assign R1C1_N83 = R1C1_Q5;
assign R1C1_S83 = R1C1_Q5;
assign R1C1_N24 = R1C1_Q4;
assign R1C1_N27 = R1C1_Q7;
assign R1C1_S24 = R1C1_Q4;
assign R1C1_S27 = R1C1_Q7;
assign R1C1_N20 = R1C1_Q0;
assign R1C1_N23 = R1C1_Q3;
assign R1C1_S20 = R1C1_Q0;
assign R1C1_S23 = R1C1_Q3;
assign R1C1_N80 = R1C1_Q0;
assign R1C1_S80 = R1C1_Q0;
assign R1C1_E83 = R1C1_Q5;
assign R1C1_W83 = R1C1_Q5;
assign R1C1_E25 = R1C1_Q5;
assign R1C1_E26 = R1C1_Q6;
assign R1C1_W25 = R1C1_Q5;
assign R1C1_W26 = R1C1_Q6;
assign R1C1_E24 = R1C1_Q4;
assign R1C1_E27 = R1C1_Q7;
assign R1C1_W24 = R1C1_Q4;
assign R1C1_W27 = R1C1_Q7;
assign R1C1_E20 = R1C1_Q0;
assign R1C1_E23 = R1C1_Q3;
assign R1C1_W20 = R1C1_Q0;
assign R1C1_W23 = R1C1_Q3;
assign R1C1_B0 = R1C1_F3;
assign R1C1_B1 = R1C1_F3;
assign R1C1_B2 = R1C1_F1;
assign R1C1_B3 = R1C1_F1;
assign R1C1_B4 = R1C1_F1;
assign R1C1_B5 = R1C1_F1;
assign R1C1_B6 = R1C1_F1;
assign R1C1_B7 = R1C1_F1;
assign R1C1_D0 = R1C1_F2;
assign R1C1_D1 = R1C1_F2;
assign R1C1_D2 = R1C1_F0;
assign R1C1_D3 = R1C1_F0;
assign R1C1_D4 = R1C1_F0;
assign R1C1_D5 = R1C1_F0;
assign R1C1_D6 = R1C1_F0;
assign R1C1_D7 = R1C1_F0;
assign R1C1_X02 = R1C1_Q1;
assign R1C1_X04 = R1C1_Q7;
assign R1C1_X06 = R1C1_Q1;
assign R1C1_X08 = R1C1_Q7;
assign R1C1_X01 = R1C1_Q0;
assign R1C1_X03 = R1C1_Q6;
assign R1C1_X05 = R1C1_Q0;
assign R1C1_X07 = R1C1_Q6;
assign R1C1_N10 = R1C1_Q0;
assign R1C1_SN10 = R1C1_Q0;
assign R1C1_SN20 = R1C1_Q0;
assign R1C1_N13 = R1C1_Q0;
assign R1C1_S10 = R1C1_Q0;
assign R1C1_S13 = R1C1_Q0;
assign R1C1_E10 = R1C1_Q0;
assign R1C1_EW10 = R1C1_Q0;
assign R1C1_EW20 = R1C1_Q0;
assign R1C1_E13 = R1C1_Q0;
assign R1C1_W10 = R1C1_Q0;
assign R1C1_W13 = R1C1_Q0;
assign R1C1_E11 = R1C1_EW10;
assign R1C1_W11 = R1C1_EW10;
assign R1C1_E12 = R1C1_EW20;
assign R1C1_W12 = R1C1_EW20;
assign R1C1_S11 = R1C1_SN10;
assign R1C1_N11 = R1C1_SN10;
assign R1C1_S12 = R1C1_SN20;
assign R1C1_N12 = R1C1_SN20;
assign VCC = 1;
assign GND = 0;
assign R1C47_CLK0 = VCC;
assign R1C47_CLK1 = VCC;
assign R1C47_CLK2 = VCC;
assign R1C47_LSR0 = VCC;
assign R1C47_LSR1 = VCC;
assign R1C47_LSR2 = VCC;
assign R1C47_CE0 = VCC;
assign R1C47_CE1 = VCC;
assign R1C47_CE2 = VCC;
assign R1C47_SEL0 = VCC;
assign R1C47_SEL1 = VCC;
assign R1C47_SEL2 = VCC;
assign R1C47_SEL3 = VCC;
assign R1C47_SEL4 = VCC;
assign R1C47_SEL5 = VCC;
assign R1C47_SEL6 = VCC;
assign R1C47_SEL7 = VCC;
assign R1C47_C0 = R1C47_F4;
assign R1C47_C1 = R1C47_F4;
assign R1C47_C2 = R1C47_F4;
assign R1C47_C3 = R1C47_F4;
assign R1C47_A4 = R1C47_F7;
assign R1C47_A5 = R1C47_F7;
assign R1C47_A6 = R1C47_F5;
assign R1C47_A7 = R1C47_F5;
assign R1C47_N82 = R1C47_Q4;
assign R1C47_S82 = R1C47_Q4;
assign R1C47_E82 = R1C47_Q4;
assign R1C47_W82 = R1C47_Q4;
assign R1C47_A0 = R1C47_F5;
assign R1C47_A1 = R1C47_F5;
assign R1C47_A2 = R1C47_F5;
assign R1C47_A3 = R1C47_F5;
assign R1C47_C4 = R1C47_F6;
assign R1C47_C5 = R1C47_F6;
assign R1C47_C6 = R1C47_F4;
assign R1C47_C7 = R1C47_F4;
assign R1C47_N81 = R1C47_Q1;
assign R1C47_S81 = R1C47_Q1;
assign R1C47_E81 = R1C47_Q1;
assign R1C47_W81 = R1C47_Q1;
assign R1C47_N21 = R1C47_Q1;
assign R1C47_N22 = R1C47_Q2;
assign R1C47_S21 = R1C47_Q1;
assign R1C47_S22 = R1C47_Q2;
assign R1C47_E21 = R1C47_Q1;
assign R1C47_E22 = R1C47_Q2;
assign R1C47_W21 = R1C47_Q1;
assign R1C47_W22 = R1C47_Q2;
assign R1C47_E80 = R1C47_Q0;
assign R1C47_W80 = R1C47_Q0;
assign R1C47_N25 = R1C47_Q5;
assign R1C47_N26 = R1C47_Q6;
assign R1C47_S25 = R1C47_Q5;
assign R1C47_S26 = R1C47_Q6;
assign R1C47_N83 = R1C47_Q5;
assign R1C47_S83 = R1C47_Q5;
assign R1C47_N24 = R1C47_Q4;
assign R1C47_N27 = R1C47_Q7;
assign R1C47_S24 = R1C47_Q4;
assign R1C47_S27 = R1C47_Q7;
assign R1C47_N20 = R1C47_Q0;
assign R1C47_N23 = R1C47_Q3;
assign R1C47_S20 = R1C47_Q0;
assign R1C47_S23 = R1C47_Q3;
assign R1C47_N80 = R1C47_Q0;
assign R1C47_S80 = R1C47_Q0;
assign R1C47_E83 = R1C47_Q5;
assign R1C47_W83 = R1C47_Q5;
assign R1C47_E25 = R1C47_Q5;
assign R1C47_E26 = R1C47_Q6;
assign R1C47_W25 = R1C47_Q5;
assign R1C47_W26 = R1C47_Q6;
assign R1C47_E24 = R1C47_Q4;
assign R1C47_E27 = R1C47_Q7;
assign R1C47_W24 = R1C47_Q4;
assign R1C47_W27 = R1C47_Q7;
assign R1C47_E20 = R1C47_Q0;
assign R1C47_E23 = R1C47_Q3;
assign R1C47_W20 = R1C47_Q0;
assign R1C47_W23 = R1C47_Q3;
assign R1C47_B0 = R1C47_F3;
assign R1C47_B1 = R1C47_F3;
assign R1C47_B2 = R1C47_F1;
assign R1C47_B3 = R1C47_F1;
assign R1C47_B4 = R1C47_F1;
assign R1C47_B5 = R1C47_F1;
assign R1C47_B6 = R1C47_F1;
assign R1C47_B7 = R1C47_F1;
assign R1C47_D0 = R1C47_F2;
assign R1C47_D1 = R1C47_F2;
assign R1C47_D2 = R1C47_F0;
assign R1C47_D3 = R1C47_F0;
assign R1C47_D4 = R1C47_F0;
assign R1C47_D5 = R1C47_F0;
assign R1C47_D6 = R1C47_F0;
assign R1C47_D7 = R1C47_F0;
assign R1C47_X02 = R1C47_Q1;
assign R1C47_X04 = R1C47_Q7;
assign R1C47_X06 = R1C47_Q1;
assign R1C47_X08 = R1C47_Q7;
assign R1C47_X01 = R1C47_Q0;
assign R1C47_X03 = R1C47_Q6;
assign R1C47_X05 = R1C47_Q0;
assign R1C47_X07 = R1C47_Q6;
assign R1C47_N10 = R1C47_Q0;
assign R1C47_SN10 = R1C47_Q0;
assign R1C47_SN20 = R1C47_Q0;
assign R1C47_N13 = R1C47_Q0;
assign R1C47_S10 = R1C47_Q0;
assign R1C47_S13 = R1C47_Q0;
assign R1C47_E10 = R1C47_Q0;
assign R1C47_EW10 = R1C47_Q0;
assign R1C47_EW20 = R1C47_Q0;
assign R1C47_E13 = R1C47_Q0;
assign R1C47_W10 = R1C47_Q0;
assign R1C47_W13 = R1C47_Q0;
assign R1C47_E11 = R1C47_EW10;
assign R1C47_W11 = R1C47_EW10;
assign R1C47_E12 = R1C47_EW20;
assign R1C47_W12 = R1C47_EW20;
assign R1C47_S11 = R1C47_SN10;
assign R1C47_N11 = R1C47_SN10;
assign R1C47_S12 = R1C47_SN20;
assign R1C47_N12 = R1C47_SN20;
assign R1C28_CLK0 = VCC;
assign R1C28_CLK1 = VCC;
assign R1C28_CLK2 = VCC;
assign R1C28_LSR0 = VCC;
assign R1C28_LSR1 = VCC;
assign R1C28_LSR2 = VCC;
assign R1C28_CE0 = VCC;
assign R1C28_CE1 = VCC;
assign R1C28_CE2 = VCC;
assign R1C28_SEL0 = VCC;
assign R1C28_SEL1 = VCC;
assign R1C28_SEL2 = VCC;
assign R1C28_SEL3 = VCC;
assign R1C28_SEL4 = VCC;
assign R1C28_SEL5 = VCC;
assign R1C28_SEL6 = VCC;
assign R1C28_SEL7 = VCC;
assign R1C28_C0 = R1C28_F4;
assign R1C28_C1 = R1C28_F4;
assign R1C28_C2 = R1C28_F4;
assign R1C28_C3 = R1C28_F4;
assign R1C28_A4 = R1C28_F7;
assign R1C28_A5 = R1C28_F7;
assign R1C28_A6 = R1C28_F5;
assign R1C28_A7 = R1C28_F5;
assign R1C28_N82 = R1C28_Q4;
assign R1C28_S82 = R1C28_Q4;
assign R1C28_E82 = R1C28_Q4;
assign R1C28_W82 = R1C28_Q4;
assign R1C28_A0 = R1C28_F5;
assign R1C28_A1 = R1C28_F5;
assign R1C28_A2 = R1C28_F5;
assign R1C28_A3 = R1C28_F5;
assign R1C28_C4 = R1C28_F6;
assign R1C28_C5 = R1C28_F6;
assign R1C28_C6 = R1C28_F4;
assign R1C28_C7 = R1C28_F4;
assign R1C28_N81 = R1C28_Q1;
assign R1C28_S81 = R1C28_Q1;
assign R1C28_E81 = R1C28_Q1;
assign R1C28_W81 = R1C28_Q1;
assign R1C28_N21 = R1C28_Q1;
assign R1C28_N22 = R1C28_Q2;
assign R1C28_S21 = R1C28_Q1;
assign R1C28_S22 = R1C28_Q2;
assign R1C28_E21 = R1C28_Q1;
assign R1C28_E22 = R1C28_Q2;
assign R1C28_W21 = R1C28_Q1;
assign R1C28_W22 = R1C28_Q2;
assign R1C28_E80 = R1C28_Q0;
assign R1C28_W80 = R1C28_Q0;
assign R1C28_N25 = R1C28_Q5;
assign R1C28_N26 = R1C28_Q6;
assign R1C28_S25 = R1C28_Q5;
assign R1C28_S26 = R1C28_Q6;
assign R1C28_N83 = R1C28_Q5;
assign R1C28_S83 = R1C28_Q5;
assign R1C28_N24 = R1C28_Q4;
assign R1C28_N27 = R1C28_Q7;
assign R1C28_S24 = R1C28_Q4;
assign R1C28_S27 = R1C28_Q7;
assign R1C28_N20 = R1C28_Q0;
assign R1C28_N23 = R1C28_Q3;
assign R1C28_S20 = R1C28_Q0;
assign R1C28_S23 = R1C28_Q3;
assign R1C28_N80 = R1C28_Q0;
assign R1C28_S80 = R1C28_Q0;
assign R1C28_E83 = R1C28_Q5;
assign R1C28_W83 = R1C28_Q5;
assign R1C28_E25 = R1C28_Q5;
assign R1C28_E26 = R1C28_Q6;
assign R1C28_W25 = R1C28_Q5;
assign R1C28_W26 = R1C28_Q6;
assign R1C28_E24 = R1C28_Q4;
assign R1C28_E27 = R1C28_Q7;
assign R1C28_W24 = R1C28_Q4;
assign R1C28_W27 = R1C28_Q7;
assign R1C28_E20 = R1C28_Q0;
assign R1C28_E23 = R1C28_Q3;
assign R1C28_W20 = R1C28_Q0;
assign R1C28_W23 = R1C28_Q3;
assign R1C28_B0 = R1C28_F3;
assign R1C28_B1 = R1C28_F3;
assign R1C28_B2 = R1C28_F1;
assign R1C28_B3 = R1C28_F1;
assign R1C28_B4 = R1C28_F1;
assign R1C28_B5 = R1C28_F1;
assign R1C28_B6 = R1C28_F1;
assign R1C28_B7 = R1C28_F1;
assign R1C28_D0 = R1C28_F2;
assign R1C28_D1 = R1C28_F2;
assign R1C28_D2 = R1C28_F0;
assign R1C28_D3 = R1C28_F0;
assign R1C28_D4 = R1C28_F0;
assign R1C28_D5 = R1C28_F0;
assign R1C28_D6 = R1C28_F0;
assign R1C28_D7 = R1C28_F0;
assign R1C28_X02 = R1C28_Q1;
assign R1C28_X04 = R1C28_Q7;
assign R1C28_X06 = R1C28_Q1;
assign R1C28_X08 = R1C28_Q7;
assign R1C28_X01 = R1C28_Q0;
assign R1C28_X03 = R1C28_Q6;
assign R1C28_X05 = R1C28_Q0;
assign R1C28_X07 = R1C28_Q6;
assign R1C28_N10 = R1C28_Q0;
assign R1C28_SN10 = R1C28_Q0;
assign R1C28_SN20 = R1C28_Q0;
assign R1C28_N13 = R1C28_Q0;
assign R1C28_S10 = R1C28_Q0;
assign R1C28_S13 = R1C28_Q0;
assign R1C28_E10 = R1C28_Q0;
assign R1C28_EW10 = R1C28_Q0;
assign R1C28_EW20 = R1C28_Q0;
assign R1C28_E13 = R1C28_Q0;
assign R1C28_W10 = R1C28_Q0;
assign R1C28_W13 = R1C28_Q0;
assign R1C28_E11 = R1C28_EW10;
assign R1C28_W11 = R1C28_EW10;
assign R1C28_E12 = R1C28_EW20;
assign R1C28_W12 = R1C28_EW20;
assign R1C28_S11 = R1C28_SN10;
assign R1C28_N11 = R1C28_SN10;
assign R1C28_S12 = R1C28_SN20;
assign R1C28_N12 = R1C28_SN20;
assign R1C32_CLK0 = VCC;
assign R1C32_CLK1 = VCC;
assign R1C32_CLK2 = VCC;
assign R1C32_LSR0 = VCC;
assign R1C32_LSR1 = VCC;
assign R1C32_LSR2 = VCC;
assign R1C32_CE0 = VCC;
assign R1C32_CE1 = VCC;
assign R1C32_CE2 = VCC;
assign R1C32_SEL0 = VCC;
assign R1C32_SEL1 = VCC;
assign R1C32_SEL2 = VCC;
assign R1C32_SEL3 = VCC;
assign R1C32_SEL4 = VCC;
assign R1C32_SEL5 = VCC;
assign R1C32_SEL6 = VCC;
assign R1C32_SEL7 = VCC;
assign R1C32_C0 = R1C32_F4;
assign R1C32_C1 = R1C32_F4;
assign R1C32_C2 = R1C32_F4;
assign R1C32_C3 = R1C32_F4;
assign R1C32_A4 = R1C32_F7;
assign R1C32_A5 = R1C32_F7;
assign R1C32_A6 = R1C32_F5;
assign R1C32_A7 = R1C32_F5;
assign R1C32_N82 = R1C32_Q4;
assign R1C32_S82 = R1C32_Q4;
assign R1C32_E82 = R1C32_Q4;
assign R1C32_W82 = R1C32_Q4;
assign R1C32_A0 = R1C32_E21;
assign R1C32_A1 = R1C32_F5;
assign R1C32_A2 = R1C32_F5;
assign R1C32_A3 = R1C32_F5;
assign R1C32_C4 = R1C32_F6;
assign R1C32_C5 = R1C32_F6;
assign R1C32_C6 = R1C32_F4;
assign R1C32_C7 = R1C32_F4;
assign R1C32_N81 = R1C32_Q1;
assign R1C32_S81 = R1C32_Q1;
assign R1C32_E81 = R1C32_Q1;
assign R1C32_W81 = R1C32_Q1;
assign R1C32_N21 = R1C32_Q1;
assign R1C32_N22 = R1C32_Q2;
assign R1C32_S21 = R1C32_Q1;
assign R1C32_S22 = R1C32_Q2;
assign R1C32_E21 = VSS;
assign R1C32_E22 = R1C32_Q2;
assign R1C32_W21 = R1C32_Q1;
assign R1C32_W22 = R1C32_Q2;
assign R1C32_E80 = R1C32_Q0;
assign R1C32_W80 = R1C32_Q0;
assign R1C32_N25 = R1C32_Q5;
assign R1C32_N26 = R1C32_Q6;
assign R1C32_S25 = R1C32_Q5;
assign R1C32_S26 = R1C32_Q6;
assign R1C32_N83 = R1C32_Q5;
assign R1C32_S83 = R1C32_Q5;
assign R1C32_N24 = R1C32_Q4;
assign R1C32_N27 = R1C32_Q7;
assign R1C32_S24 = VCC;
assign R1C32_S27 = R1C32_Q7;
assign R1C32_N20 = R1C32_Q0;
assign R1C32_N23 = R1C32_Q3;
assign R1C32_S20 = R1C32_Q0;
assign R1C32_S23 = R1C32_Q3;
assign R1C32_N80 = R1C32_Q0;
assign R1C32_S80 = R1C32_Q0;
assign R1C32_E83 = R1C32_Q5;
assign R1C32_W83 = R1C32_Q5;
assign R1C32_E25 = R1C32_Q5;
assign R1C32_E26 = R1C32_Q6;
assign R1C32_W25 = R1C32_Q5;
assign R1C32_W26 = R1C32_Q6;
assign R1C32_E24 = R1C32_Q4;
assign R1C32_E27 = R1C32_Q7;
assign R1C32_W24 = R1C32_Q4;
assign R1C32_W27 = R1C32_Q7;
assign R1C32_E20 = R1C32_Q0;
assign R1C32_E23 = R1C32_Q3;
assign R1C32_W20 = R1C32_Q0;
assign R1C32_W23 = R1C32_Q3;
assign R1C32_B0 = R1C32_S24;
assign R1C32_B1 = R1C32_F3;
assign R1C32_B2 = R1C32_F1;
assign R1C32_B3 = R1C32_F1;
assign R1C32_B4 = R1C32_F1;
assign R1C32_B5 = R1C32_F1;
assign R1C32_B6 = R1C32_F1;
assign R1C32_B7 = R1C32_F1;
assign R1C32_D0 = R1C32_F2;
assign R1C32_D1 = R1C32_F2;
assign R1C32_D2 = R1C32_F0;
assign R1C32_D3 = R1C32_F0;
assign R1C32_D4 = R1C32_F0;
assign R1C32_D5 = R1C32_F0;
assign R1C32_D6 = R1C32_F0;
assign R1C32_D7 = R1C32_F0;
assign R1C32_X02 = R1C32_Q1;
assign R1C32_X04 = R1C32_Q7;
assign R1C32_X06 = R1C32_Q1;
assign R1C32_X08 = R1C32_Q7;
assign R1C32_X01 = R1C32_Q0;
assign R1C32_X03 = R1C32_Q6;
assign R1C32_X05 = R1C32_Q0;
assign R1C32_X07 = R1C32_Q6;
assign R1C32_N10 = R1C32_Q0;
assign R1C32_SN10 = R1C32_Q0;
assign R1C32_SN20 = R1C32_Q0;
assign R1C32_N13 = R1C32_Q0;
assign R1C32_S10 = R1C32_Q0;
assign R1C32_S13 = R1C32_Q0;
assign R1C32_E10 = R1C32_Q0;
assign R1C32_EW10 = R1C32_Q0;
assign R1C32_EW20 = R1C32_Q0;
assign R1C32_E13 = R1C32_Q0;
assign R1C32_W10 = R1C32_Q0;
assign R1C32_W13 = R1C32_Q0;
assign R1C32_E11 = R1C32_EW10;
assign R1C32_W11 = R1C32_EW10;
assign R1C32_E12 = R1C32_EW20;
assign R1C32_W12 = R1C32_EW20;
assign R1C32_S11 = R1C32_SN10;
assign R1C32_N11 = R1C32_SN10;
assign R1C32_S12 = R1C32_SN20;
assign R1C32_N12 = R1C32_SN20;
assign R10C7_CLK0 = VCC;
assign R10C7_CLK1 = VCC;
assign R10C7_CLK2 = VCC;
assign R10C7_LSR0 = VCC;
assign R10C7_LSR1 = VCC;
assign R10C7_LSR2 = VCC;
assign R10C7_CE0 = VCC;
assign R10C7_CE1 = VCC;
assign R10C7_CE2 = VCC;
assign R10C7_SEL0 = VCC;
assign R10C7_SEL1 = VCC;
assign R10C7_SEL2 = VCC;
assign R10C7_SEL3 = VCC;
assign R10C7_SEL4 = VCC;
assign R10C7_SEL5 = VCC;
assign R10C7_SEL6 = VCC;
assign R10C7_SEL7 = VCC;
assign R10C7_C0 = R10C7_F4;
assign R10C7_C1 = R10C7_F4;
assign R10C7_C2 = R10C7_F4;
assign R10C7_C3 = R10C7_F4;
assign R10C7_A4 = R10C7_F7;
assign R10C7_A5 = R10C7_F7;
assign R10C7_A6 = R10C7_F5;
assign R10C7_A7 = R10C7_F5;
assign R10C7_N82 = R10C7_Q4;
assign R10C7_S82 = R10C7_Q4;
assign R10C7_E82 = R10C7_Q4;
assign R10C7_W82 = R10C7_Q4;
assign R10C7_A0 = R10C7_F5;
assign R10C7_A1 = R10C7_F5;
assign R10C7_A2 = R10C7_F5;
assign R10C7_A3 = R10C7_F5;
assign R10C7_C4 = R10C7_F6;
assign R10C7_C5 = R10C7_F6;
assign R10C7_C6 = R10C7_F4;
assign R10C7_C7 = R10C7_F4;
assign R10C7_N81 = R10C7_Q1;
assign R10C7_S81 = R10C7_Q1;
assign R10C7_E81 = R10C7_Q1;
assign R10C7_W81 = R10C7_Q1;
assign R10C7_N21 = R10C7_Q1;
assign R10C7_N22 = R10C7_Q2;
assign R10C7_S21 = R10C7_Q1;
assign R10C7_S22 = R10C7_Q2;
assign R10C7_E21 = R10C7_Q1;
assign R10C7_E22 = R10C7_Q2;
assign R10C7_W21 = R10C7_Q1;
assign R10C7_W22 = R10C7_Q2;
assign R10C7_E80 = R10C7_Q0;
assign R10C7_W80 = R10C7_Q0;
assign R10C7_N25 = R10C7_Q5;
assign R10C7_N26 = R10C7_Q6;
assign R10C7_S25 = R10C7_Q5;
assign R10C7_S26 = R10C7_Q6;
assign R10C7_N83 = R10C7_Q5;
assign R10C7_S83 = R10C7_Q5;
assign R10C7_N24 = R10C7_Q4;
assign R10C7_N27 = R10C7_Q7;
assign R10C7_S24 = R10C7_Q4;
assign R10C7_S27 = R10C7_Q7;
assign R10C7_N20 = R10C7_Q0;
assign R10C7_N23 = R10C7_Q3;
assign R10C7_S20 = R10C7_Q0;
assign R10C7_S23 = R10C7_Q3;
assign R10C7_N80 = R10C7_Q0;
assign R10C7_S80 = R10C7_Q0;
assign R10C7_E83 = R10C7_Q5;
assign R10C7_W83 = R10C7_Q5;
assign R10C7_E25 = R10C7_Q5;
assign R10C7_E26 = R10C7_Q6;
assign R10C7_W25 = R10C7_Q5;
assign R10C7_W26 = R10C7_Q6;
assign R10C7_E24 = R10C7_Q4;
assign R10C7_E27 = R10C7_Q7;
assign R10C7_W24 = R10C7_Q4;
assign R10C7_W27 = R10C7_Q7;
assign R10C7_E20 = R10C7_Q0;
assign R10C7_E23 = R10C7_Q3;
assign R10C7_W20 = R10C7_Q0;
assign R10C7_W23 = R10C7_Q3;
assign R10C7_B0 = R10C7_F3;
assign R10C7_B1 = R10C7_F3;
assign R10C7_B2 = R10C7_F1;
assign R10C7_B3 = R10C7_F1;
assign R10C7_B4 = R10C7_F1;
assign R10C7_B5 = R10C7_F1;
assign R10C7_B6 = R10C7_F1;
assign R10C7_B7 = R10C7_F1;
assign R10C7_D0 = R10C7_F2;
assign R10C7_D1 = R10C7_F2;
assign R10C7_D2 = R10C7_F0;
assign R10C7_D3 = R10C7_F0;
assign R10C7_D4 = R10C7_F0;
assign R10C7_D5 = R10C7_F0;
assign R10C7_D6 = R10C7_F0;
assign R10C7_D7 = R10C7_F0;
assign R10C7_X02 = R10C7_Q1;
assign R10C7_X04 = R10C7_Q7;
assign R10C7_X06 = R10C7_Q1;
assign R10C7_X08 = R10C7_Q7;
assign R10C7_X01 = R10C7_Q0;
assign R10C7_X03 = R10C7_Q6;
assign R10C7_X05 = R10C7_Q0;
assign R10C7_X07 = R10C7_Q6;
assign R10C7_N10 = R10C7_Q0;
assign R10C7_SN10 = R10C7_Q0;
assign R10C7_SN20 = R10C7_Q0;
assign R10C7_N13 = R10C7_Q0;
assign R10C7_S10 = R10C7_Q0;
assign R10C7_S13 = R10C7_Q0;
assign R10C7_E10 = R10C7_Q0;
assign R10C7_EW10 = R10C7_Q0;
assign R10C7_EW20 = R10C7_Q0;
assign R10C7_E13 = R10C7_Q0;
assign R10C7_W10 = R10C7_Q0;
assign R10C7_W13 = R10C7_Q0;
assign R10C7_E11 = R10C7_EW10;
assign R10C7_W11 = R10C7_EW10;
assign R10C7_E12 = R10C7_EW20;
assign R10C7_W12 = R10C7_EW20;
assign R10C7_S11 = R10C7_SN10;
assign R10C7_N11 = R10C7_SN10;
assign R10C7_S12 = R10C7_SN20;
assign R10C7_N12 = R10C7_SN20;
assign R10C10_CLK0 = VCC;
assign R10C10_CLK1 = VCC;
assign R10C10_CLK2 = VCC;
assign R10C10_LSR0 = VCC;
assign R10C10_LSR1 = VCC;
assign R10C10_LSR2 = VCC;
assign R10C10_CE0 = VCC;
assign R10C10_CE1 = VCC;
assign R10C10_CE2 = VCC;
assign R10C10_SEL0 = VCC;
assign R10C10_SEL1 = VCC;
assign R10C10_SEL2 = VCC;
assign R10C10_SEL3 = VCC;
assign R10C10_SEL4 = VCC;
assign R10C10_SEL5 = VCC;
assign R10C10_SEL6 = VCC;
assign R10C10_SEL7 = VCC;
assign R10C10_C0 = R10C10_F4;
assign R10C10_C1 = R10C10_F4;
assign R10C10_C2 = R10C10_F4;
assign R10C10_C3 = R10C10_F4;
assign R10C10_A4 = R10C10_F7;
assign R10C10_A5 = R10C10_F7;
assign R10C10_A6 = R10C10_F5;
assign R10C10_A7 = R10C10_F5;
assign R10C10_N82 = R10C10_Q4;
assign R10C10_S82 = R10C10_Q4;
assign R10C10_E82 = R10C10_Q4;
assign R10C10_W82 = R10C10_Q4;
assign R10C10_A0 = R10C10_F5;
assign R10C10_A1 = R10C10_F5;
assign R10C10_A2 = R10C10_F5;
assign R10C10_A3 = R10C10_F5;
assign R10C10_C4 = R10C10_F6;
assign R10C10_C5 = R10C10_F6;
assign R10C10_C6 = R10C10_F4;
assign R10C10_C7 = R10C10_F4;
assign R10C10_N81 = R10C10_Q1;
assign R10C10_S81 = R10C10_Q1;
assign R10C10_E81 = R10C10_Q1;
assign R10C10_W81 = R10C10_Q1;
assign R10C10_N21 = R10C10_Q1;
assign R10C10_N22 = R10C10_Q2;
assign R10C10_S21 = R10C10_Q1;
assign R10C10_S22 = R10C10_Q2;
assign R10C10_E21 = R10C10_Q1;
assign R10C10_E22 = R10C10_Q2;
assign R10C10_W21 = R10C10_Q1;
assign R10C10_W22 = R10C10_Q2;
assign R10C10_E80 = R10C10_Q0;
assign R10C10_W80 = R10C10_Q0;
assign R10C10_N25 = R10C10_Q5;
assign R10C10_N26 = R10C10_Q6;
assign R10C10_S25 = R10C10_Q5;
assign R10C10_S26 = R10C10_Q6;
assign R10C10_N83 = R10C10_Q5;
assign R10C10_S83 = R10C10_Q5;
assign R10C10_N24 = R10C10_Q4;
assign R10C10_N27 = R10C10_Q7;
assign R10C10_S24 = R10C10_Q4;
assign R10C10_S27 = R10C10_Q7;
assign R10C10_N20 = R10C10_Q0;
assign R10C10_N23 = R10C10_Q3;
assign R10C10_S20 = R10C10_Q0;
assign R10C10_S23 = R10C10_Q3;
assign R10C10_N80 = R10C10_Q0;
assign R10C10_S80 = R10C10_Q0;
assign R10C10_E83 = R10C10_Q5;
assign R10C10_W83 = R10C10_Q5;
assign R10C10_E25 = R10C10_Q5;
assign R10C10_E26 = R10C10_Q6;
assign R10C10_W25 = R10C10_Q5;
assign R10C10_W26 = R10C10_Q6;
assign R10C10_E24 = R10C10_Q4;
assign R10C10_E27 = R10C10_Q7;
assign R10C10_W24 = R10C10_Q4;
assign R10C10_W27 = R10C10_Q7;
assign R10C10_E20 = R10C10_Q0;
assign R10C10_E23 = R10C10_Q3;
assign R10C10_W20 = R10C10_Q0;
assign R10C10_W23 = R10C10_Q3;
assign R10C10_B0 = R10C10_F3;
assign R10C10_B1 = R10C10_F3;
assign R10C10_B2 = R10C10_F1;
assign R10C10_B3 = R10C10_F1;
assign R10C10_B4 = R10C10_F1;
assign R10C10_B5 = R10C10_F1;
assign R10C10_B6 = R10C10_F1;
assign R10C10_B7 = R10C10_F1;
assign R10C10_D0 = R10C10_F2;
assign R10C10_D1 = R10C10_F2;
assign R10C10_D2 = R10C10_F0;
assign R10C10_D3 = R10C10_F0;
assign R10C10_D4 = R10C10_F0;
assign R10C10_D5 = R10C10_F0;
assign R10C10_D6 = R10C10_F0;
assign R10C10_D7 = R10C10_F0;
assign R10C10_X02 = R10C10_Q1;
assign R10C10_X04 = R10C10_Q7;
assign R10C10_X06 = R10C10_Q1;
assign R10C10_X08 = R10C10_Q7;
assign R10C10_X01 = R10C10_Q0;
assign R10C10_X03 = R10C10_Q6;
assign R10C10_X05 = R10C10_Q0;
assign R10C10_X07 = R10C10_Q6;
assign R10C10_N10 = R10C10_Q0;
assign R10C10_SN10 = R10C10_Q0;
assign R10C10_SN20 = R10C10_Q0;
assign R10C10_N13 = R10C10_Q0;
assign R10C10_S10 = R10C10_Q0;
assign R10C10_S13 = R10C10_Q0;
assign R10C10_E10 = R10C10_Q0;
assign R10C10_EW10 = R10C10_Q0;
assign R10C10_EW20 = R10C10_Q0;
assign R10C10_E13 = R10C10_Q0;
assign R10C10_W10 = R10C10_Q0;
assign R10C10_W13 = R10C10_Q0;
assign R10C10_E11 = R10C10_EW10;
assign R10C10_W11 = R10C10_EW10;
assign R10C10_E12 = R10C10_EW20;
assign R10C10_W12 = R10C10_EW20;
assign R10C10_S11 = R10C10_SN10;
assign R10C10_N11 = R10C10_SN10;
assign R10C10_S12 = R10C10_SN20;
assign R10C10_N12 = R10C10_SN20;
assign R10C13_CLK0 = VCC;
assign R10C13_CLK1 = VCC;
assign R10C13_CLK2 = VCC;
assign R10C13_LSR0 = VCC;
assign R10C13_LSR1 = VCC;
assign R10C13_LSR2 = VCC;
assign R10C13_CE0 = VCC;
assign R10C13_CE1 = VCC;
assign R10C13_CE2 = VCC;
assign R10C13_SEL0 = VCC;
assign R10C13_SEL1 = VCC;
assign R10C13_SEL2 = VCC;
assign R10C13_SEL3 = VCC;
assign R10C13_SEL4 = VCC;
assign R10C13_SEL5 = VCC;
assign R10C13_SEL6 = VCC;
assign R10C13_SEL7 = VCC;
assign R10C13_C0 = R10C13_F4;
assign R10C13_C1 = R10C13_F4;
assign R10C13_C2 = R10C13_F4;
assign R10C13_C3 = R10C13_F4;
assign R10C13_A4 = R10C13_F7;
assign R10C13_A5 = R10C13_F7;
assign R10C13_A6 = R10C13_F5;
assign R10C13_A7 = R10C13_F5;
assign R10C13_N82 = R10C13_Q4;
assign R10C13_S82 = R10C13_Q4;
assign R10C13_E82 = R10C13_Q4;
assign R10C13_W82 = R10C13_Q4;
assign R10C13_A0 = R10C13_F5;
assign R10C13_A1 = R10C13_F5;
assign R10C13_A2 = R10C13_F5;
assign R10C13_A3 = R10C13_F5;
assign R10C13_C4 = R10C13_F6;
assign R10C13_C5 = R10C13_F6;
assign R10C13_C6 = R10C13_F4;
assign R10C13_C7 = R10C13_F4;
assign R10C13_N81 = R10C13_Q1;
assign R10C13_S81 = R10C13_Q1;
assign R10C13_E81 = R10C13_Q1;
assign R10C13_W81 = R10C13_Q1;
assign R10C13_N21 = R10C13_Q1;
assign R10C13_N22 = R10C13_Q2;
assign R10C13_S21 = R10C13_Q1;
assign R10C13_S22 = R10C13_Q2;
assign R10C13_E21 = R10C13_Q1;
assign R10C13_E22 = R10C13_Q2;
assign R10C13_W21 = R10C13_Q1;
assign R10C13_W22 = R10C13_Q2;
assign R10C13_E80 = R10C13_Q0;
assign R10C13_W80 = R10C13_Q0;
assign R10C13_N25 = R10C13_Q5;
assign R10C13_N26 = R10C13_Q6;
assign R10C13_S25 = R10C13_Q5;
assign R10C13_S26 = R10C13_Q6;
assign R10C13_N83 = R10C13_Q5;
assign R10C13_S83 = R10C13_Q5;
assign R10C13_N24 = R10C13_Q4;
assign R10C13_N27 = R10C13_Q7;
assign R10C13_S24 = R10C13_Q4;
assign R10C13_S27 = R10C13_Q7;
assign R10C13_N20 = R10C13_Q0;
assign R10C13_N23 = R10C13_Q3;
assign R10C13_S20 = R10C13_Q0;
assign R10C13_S23 = R10C13_Q3;
assign R10C13_N80 = R10C13_Q0;
assign R10C13_S80 = R10C13_Q0;
assign R10C13_E83 = R10C13_Q5;
assign R10C13_W83 = R10C13_Q5;
assign R10C13_E25 = R10C13_Q5;
assign R10C13_E26 = R10C13_Q6;
assign R10C13_W25 = R10C13_Q5;
assign R10C13_W26 = R10C13_Q6;
assign R10C13_E24 = R10C13_Q4;
assign R10C13_E27 = R10C13_Q7;
assign R10C13_W24 = R10C13_Q4;
assign R10C13_W27 = R10C13_Q7;
assign R10C13_E20 = R10C13_Q0;
assign R10C13_E23 = R10C13_Q3;
assign R10C13_W20 = R10C13_Q0;
assign R10C13_W23 = R10C13_Q3;
assign R10C13_B0 = R10C13_F3;
assign R10C13_B1 = R10C13_F3;
assign R10C13_B2 = R10C13_F1;
assign R10C13_B3 = R10C13_F1;
assign R10C13_B4 = R10C13_F1;
assign R10C13_B5 = R10C13_F1;
assign R10C13_B6 = R10C13_F1;
assign R10C13_B7 = R10C13_F1;
assign R10C13_D0 = R10C13_F2;
assign R10C13_D1 = R10C13_F2;
assign R10C13_D2 = R10C13_F0;
assign R10C13_D3 = R10C13_F0;
assign R10C13_D4 = R10C13_F0;
assign R10C13_D5 = R10C13_F0;
assign R10C13_D6 = R10C13_F0;
assign R10C13_D7 = R10C13_F0;
assign R10C13_X02 = R10C13_Q1;
assign R10C13_X04 = R10C13_Q7;
assign R10C13_X06 = R10C13_Q1;
assign R10C13_X08 = R10C13_Q7;
assign R10C13_X01 = R10C13_Q0;
assign R10C13_X03 = R10C13_Q6;
assign R10C13_X05 = R10C13_Q0;
assign R10C13_X07 = R10C13_Q6;
assign R10C13_N10 = R10C13_Q0;
assign R10C13_SN10 = R10C13_Q0;
assign R10C13_SN20 = R10C13_Q0;
assign R10C13_N13 = R10C13_Q0;
assign R10C13_S10 = R10C13_Q0;
assign R10C13_S13 = R10C13_Q0;
assign R10C13_E10 = R10C13_Q0;
assign R10C13_EW10 = R10C13_Q0;
assign R10C13_EW20 = R10C13_Q0;
assign R10C13_E13 = R10C13_Q0;
assign R10C13_W10 = R10C13_Q0;
assign R10C13_W13 = R10C13_Q0;
assign R10C13_E11 = R10C13_EW10;
assign R10C13_W11 = R10C13_EW10;
assign R10C13_E12 = R10C13_EW20;
assign R10C13_W12 = R10C13_EW20;
assign R10C13_S11 = R10C13_SN10;
assign R10C13_N11 = R10C13_SN10;
assign R10C13_S12 = R10C13_SN20;
assign R10C13_N12 = R10C13_SN20;
assign R10C16_CLK0 = VCC;
assign R10C16_CLK1 = VCC;
assign R10C16_CLK2 = VCC;
assign R10C16_LSR0 = VCC;
assign R10C16_LSR1 = VCC;
assign R10C16_LSR2 = VCC;
assign R10C16_CE0 = VCC;
assign R10C16_CE1 = VCC;
assign R10C16_CE2 = VCC;
assign R10C16_SEL0 = VCC;
assign R10C16_SEL1 = VCC;
assign R10C16_SEL2 = VCC;
assign R10C16_SEL3 = VCC;
assign R10C16_SEL4 = VCC;
assign R10C16_SEL5 = VCC;
assign R10C16_SEL6 = VCC;
assign R10C16_SEL7 = VCC;
assign R10C16_C0 = R10C16_F4;
assign R10C16_C1 = R10C16_F4;
assign R10C16_C2 = R10C16_F4;
assign R10C16_C3 = R10C16_F4;
assign R10C16_A4 = R10C16_F7;
assign R10C16_A5 = R10C16_F7;
assign R10C16_A6 = R10C16_F5;
assign R10C16_A7 = R10C16_F5;
assign R10C16_N82 = R10C16_Q4;
assign R10C16_S82 = R10C16_Q4;
assign R10C16_E82 = R10C16_Q4;
assign R10C16_W82 = R10C16_Q4;
assign R10C16_A0 = R10C16_F5;
assign R10C16_A1 = R10C16_F5;
assign R10C16_A2 = R10C16_F5;
assign R10C16_A3 = R10C16_F5;
assign R10C16_C4 = R10C16_F6;
assign R10C16_C5 = R10C16_F6;
assign R10C16_C6 = R10C16_F4;
assign R10C16_C7 = R10C16_F4;
assign R10C16_N81 = R10C16_Q1;
assign R10C16_S81 = R10C16_Q1;
assign R10C16_E81 = R10C16_Q1;
assign R10C16_W81 = R10C16_Q1;
assign R10C16_N21 = R10C16_Q1;
assign R10C16_N22 = R10C16_Q2;
assign R10C16_S21 = R10C16_Q1;
assign R10C16_S22 = R10C16_Q2;
assign R10C16_E21 = R10C16_Q1;
assign R10C16_E22 = R10C16_Q2;
assign R10C16_W21 = R10C16_Q1;
assign R10C16_W22 = R10C16_Q2;
assign R10C16_E80 = R10C16_Q0;
assign R10C16_W80 = R10C16_Q0;
assign R10C16_N25 = R10C16_Q5;
assign R10C16_N26 = R10C16_Q6;
assign R10C16_S25 = R10C16_Q5;
assign R10C16_S26 = R10C16_Q6;
assign R10C16_N83 = R10C16_Q5;
assign R10C16_S83 = R10C16_Q5;
assign R10C16_N24 = R10C16_Q4;
assign R10C16_N27 = R10C16_Q7;
assign R10C16_S24 = R10C16_Q4;
assign R10C16_S27 = R10C16_Q7;
assign R10C16_N20 = R10C16_Q0;
assign R10C16_N23 = R10C16_Q3;
assign R10C16_S20 = R10C16_Q0;
assign R10C16_S23 = R10C16_Q3;
assign R10C16_N80 = R10C16_Q0;
assign R10C16_S80 = R10C16_Q0;
assign R10C16_E83 = R10C16_Q5;
assign R10C16_W83 = R10C16_Q5;
assign R10C16_E25 = R10C16_Q5;
assign R10C16_E26 = R10C16_Q6;
assign R10C16_W25 = R10C16_Q5;
assign R10C16_W26 = R10C16_Q6;
assign R10C16_E24 = R10C16_Q4;
assign R10C16_E27 = R10C16_Q7;
assign R10C16_W24 = R10C16_Q4;
assign R10C16_W27 = R10C16_Q7;
assign R10C16_E20 = R10C16_Q0;
assign R10C16_E23 = R10C16_Q3;
assign R10C16_W20 = R10C16_Q0;
assign R10C16_W23 = R10C16_Q3;
assign R10C16_B0 = R10C16_F3;
assign R10C16_B1 = R10C16_F3;
assign R10C16_B2 = R10C16_F1;
assign R10C16_B3 = R10C16_F1;
assign R10C16_B4 = R10C16_F1;
assign R10C16_B5 = R10C16_F1;
assign R10C16_B6 = R10C16_F1;
assign R10C16_B7 = R10C16_F1;
assign R10C16_D0 = R10C16_F2;
assign R10C16_D1 = R10C16_F2;
assign R10C16_D2 = R10C16_F0;
assign R10C16_D3 = R10C16_F0;
assign R10C16_D4 = R10C16_F0;
assign R10C16_D5 = R10C16_F0;
assign R10C16_D6 = R10C16_F0;
assign R10C16_D7 = R10C16_F0;
assign R10C16_X02 = R10C16_Q1;
assign R10C16_X04 = R10C16_Q7;
assign R10C16_X06 = R10C16_Q1;
assign R10C16_X08 = R10C16_Q7;
assign R10C16_X01 = R10C16_Q0;
assign R10C16_X03 = R10C16_Q6;
assign R10C16_X05 = R10C16_Q0;
assign R10C16_X07 = R10C16_Q6;
assign R10C16_N10 = R10C16_Q0;
assign R10C16_SN10 = R10C16_Q0;
assign R10C16_SN20 = R10C16_Q0;
assign R10C16_N13 = R10C16_Q0;
assign R10C16_S10 = R10C16_Q0;
assign R10C16_S13 = R10C16_Q0;
assign R10C16_E10 = R10C16_Q0;
assign R10C16_EW10 = R10C16_Q0;
assign R10C16_EW20 = R10C16_Q0;
assign R10C16_E13 = R10C16_Q0;
assign R10C16_W10 = R10C16_Q0;
assign R10C16_W13 = R10C16_Q0;
assign R10C16_E11 = R10C16_EW10;
assign R10C16_W11 = R10C16_EW10;
assign R10C16_E12 = R10C16_EW20;
assign R10C16_W12 = R10C16_EW20;
assign R10C16_S11 = R10C16_SN10;
assign R10C16_N11 = R10C16_SN10;
assign R10C16_S12 = R10C16_SN20;
assign R10C16_N12 = R10C16_SN20;
assign R10C19_CLK0 = VCC;
assign R10C19_CLK1 = VCC;
assign R10C19_CLK2 = VCC;
assign R10C19_LSR0 = VCC;
assign R10C19_LSR1 = VCC;
assign R10C19_LSR2 = VCC;
assign R10C19_CE0 = VCC;
assign R10C19_CE1 = VCC;
assign R10C19_CE2 = VCC;
assign R10C19_SEL0 = VCC;
assign R10C19_SEL1 = VCC;
assign R10C19_SEL2 = VCC;
assign R10C19_SEL3 = VCC;
assign R10C19_SEL4 = VCC;
assign R10C19_SEL5 = VCC;
assign R10C19_SEL6 = VCC;
assign R10C19_SEL7 = VCC;
assign R10C19_C0 = R10C19_F4;
assign R10C19_C1 = R10C19_F4;
assign R10C19_C2 = R10C19_F4;
assign R10C19_C3 = R10C19_F4;
assign R10C19_A4 = R10C19_F7;
assign R10C19_A5 = R10C19_F7;
assign R10C19_A6 = R10C19_F5;
assign R10C19_A7 = R10C19_F5;
assign R10C19_N82 = R10C19_Q4;
assign R10C19_S82 = R10C19_Q4;
assign R10C19_E82 = R10C19_Q4;
assign R10C19_W82 = R10C19_Q4;
assign R10C19_A0 = R10C19_F5;
assign R10C19_A1 = R10C19_F5;
assign R10C19_A2 = R10C19_F5;
assign R10C19_A3 = R10C19_F5;
assign R10C19_C4 = R10C19_F6;
assign R10C19_C5 = R10C19_F6;
assign R10C19_C6 = R10C19_F4;
assign R10C19_C7 = R10C19_F4;
assign R10C19_N81 = R10C19_Q1;
assign R10C19_S81 = R10C19_Q1;
assign R10C19_E81 = R10C19_Q1;
assign R10C19_W81 = R10C19_Q1;
assign R10C19_N21 = R10C19_Q1;
assign R10C19_N22 = R10C19_Q2;
assign R10C19_S21 = R10C19_Q1;
assign R10C19_S22 = R10C19_Q2;
assign R10C19_E21 = R10C19_Q1;
assign R10C19_E22 = R10C19_Q2;
assign R10C19_W21 = R10C19_Q1;
assign R10C19_W22 = R10C19_Q2;
assign R10C19_E80 = R10C19_Q0;
assign R10C19_W80 = R10C19_Q0;
assign R10C19_N25 = R10C19_Q5;
assign R10C19_N26 = R10C19_Q6;
assign R10C19_S25 = R10C19_Q5;
assign R10C19_S26 = R10C19_Q6;
assign R10C19_N83 = R10C19_Q5;
assign R10C19_S83 = R10C19_Q5;
assign R10C19_N24 = R10C19_Q4;
assign R10C19_N27 = R10C19_Q7;
assign R10C19_S24 = R10C19_Q4;
assign R10C19_S27 = R10C19_Q7;
assign R10C19_N20 = R10C19_Q0;
assign R10C19_N23 = R10C19_Q3;
assign R10C19_S20 = R10C19_Q0;
assign R10C19_S23 = R10C19_Q3;
assign R10C19_N80 = R10C19_Q0;
assign R10C19_S80 = R10C19_Q0;
assign R10C19_E83 = R10C19_Q5;
assign R10C19_W83 = R10C19_Q5;
assign R10C19_E25 = R10C19_Q5;
assign R10C19_E26 = R10C19_Q6;
assign R10C19_W25 = R10C19_Q5;
assign R10C19_W26 = R10C19_Q6;
assign R10C19_E24 = R10C19_Q4;
assign R10C19_E27 = R10C19_Q7;
assign R10C19_W24 = R10C19_Q4;
assign R10C19_W27 = R10C19_Q7;
assign R10C19_E20 = R10C19_Q0;
assign R10C19_E23 = R10C19_Q3;
assign R10C19_W20 = R10C19_Q0;
assign R10C19_W23 = R10C19_Q3;
assign R10C19_B0 = R10C19_F3;
assign R10C19_B1 = R10C19_F3;
assign R10C19_B2 = R10C19_F1;
assign R10C19_B3 = R10C19_F1;
assign R10C19_B4 = R10C19_F1;
assign R10C19_B5 = R10C19_F1;
assign R10C19_B6 = R10C19_F1;
assign R10C19_B7 = R10C19_F1;
assign R10C19_D0 = R10C19_F2;
assign R10C19_D1 = R10C19_F2;
assign R10C19_D2 = R10C19_F0;
assign R10C19_D3 = R10C19_F0;
assign R10C19_D4 = R10C19_F0;
assign R10C19_D5 = R10C19_F0;
assign R10C19_D6 = R10C19_F0;
assign R10C19_D7 = R10C19_F0;
assign R10C19_X02 = R10C19_Q1;
assign R10C19_X04 = R10C19_Q7;
assign R10C19_X06 = R10C19_Q1;
assign R10C19_X08 = R10C19_Q7;
assign R10C19_X01 = R10C19_Q0;
assign R10C19_X03 = R10C19_Q6;
assign R10C19_X05 = R10C19_Q0;
assign R10C19_X07 = R10C19_Q6;
assign R10C19_N10 = R10C19_Q0;
assign R10C19_SN10 = R10C19_Q0;
assign R10C19_SN20 = R10C19_Q0;
assign R10C19_N13 = R10C19_Q0;
assign R10C19_S10 = R10C19_Q0;
assign R10C19_S13 = R10C19_Q0;
assign R10C19_E10 = R10C19_Q0;
assign R10C19_EW10 = R10C19_Q0;
assign R10C19_EW20 = R10C19_Q0;
assign R10C19_E13 = R10C19_Q0;
assign R10C19_W10 = R10C19_Q0;
assign R10C19_W13 = R10C19_Q0;
assign R10C19_E11 = R10C19_EW10;
assign R10C19_W11 = R10C19_EW10;
assign R10C19_E12 = R10C19_EW20;
assign R10C19_W12 = R10C19_EW20;
assign R10C19_S11 = R10C19_SN10;
assign R10C19_N11 = R10C19_SN10;
assign R10C19_S12 = R10C19_SN20;
assign R10C19_N12 = R10C19_SN20;
assign R10C22_CLK0 = VCC;
assign R10C22_CLK1 = VCC;
assign R10C22_CLK2 = VCC;
assign R10C22_LSR0 = VCC;
assign R10C22_LSR1 = VCC;
assign R10C22_LSR2 = VCC;
assign R10C22_CE0 = VCC;
assign R10C22_CE1 = VCC;
assign R10C22_CE2 = VCC;
assign R10C22_SEL0 = VCC;
assign R10C22_SEL1 = VCC;
assign R10C22_SEL2 = VCC;
assign R10C22_SEL3 = VCC;
assign R10C22_SEL4 = VCC;
assign R10C22_SEL5 = VCC;
assign R10C22_SEL6 = VCC;
assign R10C22_SEL7 = VCC;
assign R10C22_C0 = R10C22_F4;
assign R10C22_C1 = R10C22_F4;
assign R10C22_C2 = R10C22_F4;
assign R10C22_C3 = R10C22_F4;
assign R10C22_A4 = R10C22_F7;
assign R10C22_A5 = R10C22_F7;
assign R10C22_A6 = R10C22_F5;
assign R10C22_A7 = R10C22_F5;
assign R10C22_N82 = R10C22_Q4;
assign R10C22_S82 = R10C22_Q4;
assign R10C22_E82 = R10C22_Q4;
assign R10C22_W82 = R10C22_Q4;
assign R10C22_A0 = R10C22_F5;
assign R10C22_A1 = R10C22_F5;
assign R10C22_A2 = R10C22_F5;
assign R10C22_A3 = R10C22_F5;
assign R10C22_C4 = R10C22_F6;
assign R10C22_C5 = R10C22_F6;
assign R10C22_C6 = R10C22_F4;
assign R10C22_C7 = R10C22_F4;
assign R10C22_N81 = R10C22_Q1;
assign R10C22_S81 = R10C22_Q1;
assign R10C22_E81 = R10C22_Q1;
assign R10C22_W81 = R10C22_Q1;
assign R10C22_N21 = R10C22_Q1;
assign R10C22_N22 = R10C22_Q2;
assign R10C22_S21 = R10C22_Q1;
assign R10C22_S22 = R10C22_Q2;
assign R10C22_E21 = R10C22_Q1;
assign R10C22_E22 = R10C22_Q2;
assign R10C22_W21 = R10C22_Q1;
assign R10C22_W22 = R10C22_Q2;
assign R10C22_E80 = R10C22_Q0;
assign R10C22_W80 = R10C22_Q0;
assign R10C22_N25 = R10C22_Q5;
assign R10C22_N26 = R10C22_Q6;
assign R10C22_S25 = R10C22_Q5;
assign R10C22_S26 = R10C22_Q6;
assign R10C22_N83 = R10C22_Q5;
assign R10C22_S83 = R10C22_Q5;
assign R10C22_N24 = R10C22_Q4;
assign R10C22_N27 = R10C22_Q7;
assign R10C22_S24 = R10C22_Q4;
assign R10C22_S27 = R10C22_Q7;
assign R10C22_N20 = R10C22_Q0;
assign R10C22_N23 = R10C22_Q3;
assign R10C22_S20 = R10C22_Q0;
assign R10C22_S23 = R10C22_Q3;
assign R10C22_N80 = R10C22_Q0;
assign R10C22_S80 = R10C22_Q0;
assign R10C22_E83 = R10C22_Q5;
assign R10C22_W83 = R10C22_Q5;
assign R10C22_E25 = R10C22_Q5;
assign R10C22_E26 = R10C22_Q6;
assign R10C22_W25 = R10C22_Q5;
assign R10C22_W26 = R10C22_Q6;
assign R10C22_E24 = R10C22_Q4;
assign R10C22_E27 = R10C22_Q7;
assign R10C22_W24 = R10C22_Q4;
assign R10C22_W27 = R10C22_Q7;
assign R10C22_E20 = R10C22_Q0;
assign R10C22_E23 = R10C22_Q3;
assign R10C22_W20 = R10C22_Q0;
assign R10C22_W23 = R10C22_Q3;
assign R10C22_B0 = R10C22_F3;
assign R10C22_B1 = R10C22_F3;
assign R10C22_B2 = R10C22_F1;
assign R10C22_B3 = R10C22_F1;
assign R10C22_B4 = R10C22_F1;
assign R10C22_B5 = R10C22_F1;
assign R10C22_B6 = R10C22_F1;
assign R10C22_B7 = R10C22_F1;
assign R10C22_D0 = R10C22_F2;
assign R10C22_D1 = R10C22_F2;
assign R10C22_D2 = R10C22_F0;
assign R10C22_D3 = R10C22_F0;
assign R10C22_D4 = R10C22_F0;
assign R10C22_D5 = R10C22_F0;
assign R10C22_D6 = R10C22_F0;
assign R10C22_D7 = R10C22_F0;
assign R10C22_X02 = R10C22_Q1;
assign R10C22_X04 = R10C22_Q7;
assign R10C22_X06 = R10C22_Q1;
assign R10C22_X08 = R10C22_Q7;
assign R10C22_X01 = R10C22_Q0;
assign R10C22_X03 = R10C22_Q6;
assign R10C22_X05 = R10C22_Q0;
assign R10C22_X07 = R10C22_Q6;
assign R10C22_N10 = R10C22_Q0;
assign R10C22_SN10 = R10C22_Q0;
assign R10C22_SN20 = R10C22_Q0;
assign R10C22_N13 = R10C22_Q0;
assign R10C22_S10 = R10C22_Q0;
assign R10C22_S13 = R10C22_Q0;
assign R10C22_E10 = R10C22_Q0;
assign R10C22_EW10 = R10C22_Q0;
assign R10C22_EW20 = R10C22_Q0;
assign R10C22_E13 = R10C22_Q0;
assign R10C22_W10 = R10C22_Q0;
assign R10C22_W13 = R10C22_Q0;
assign R10C22_E11 = R10C22_EW10;
assign R10C22_W11 = R10C22_EW10;
assign R10C22_E12 = R10C22_EW20;
assign R10C22_W12 = R10C22_EW20;
assign R10C22_S11 = R10C22_SN10;
assign R10C22_N11 = R10C22_SN10;
assign R10C22_S12 = R10C22_SN20;
assign R10C22_N12 = R10C22_SN20;
assign R10C25_CLK0 = VCC;
assign R10C25_CLK1 = VCC;
assign R10C25_CLK2 = VCC;
assign R10C25_LSR0 = VCC;
assign R10C25_LSR1 = VCC;
assign R10C25_LSR2 = VCC;
assign R10C25_CE0 = VCC;
assign R10C25_CE1 = VCC;
assign R10C25_CE2 = VCC;
assign R10C25_SEL0 = VCC;
assign R10C25_SEL1 = VCC;
assign R10C25_SEL2 = VCC;
assign R10C25_SEL3 = VCC;
assign R10C25_SEL4 = VCC;
assign R10C25_SEL5 = VCC;
assign R10C25_SEL6 = VCC;
assign R10C25_SEL7 = VCC;
assign R10C25_C0 = R10C25_F4;
assign R10C25_C1 = R10C25_F4;
assign R10C25_C2 = R10C25_F4;
assign R10C25_C3 = R10C25_F4;
assign R10C25_A4 = R10C25_F7;
assign R10C25_A5 = R10C25_F7;
assign R10C25_A6 = R10C25_F5;
assign R10C25_A7 = R10C25_F5;
assign R10C25_N82 = R10C25_Q4;
assign R10C25_S82 = R10C25_Q4;
assign R10C25_E82 = R10C25_Q4;
assign R10C25_W82 = R10C25_Q4;
assign R10C25_A0 = R10C25_F5;
assign R10C25_A1 = R10C25_F5;
assign R10C25_A2 = R10C25_F5;
assign R10C25_A3 = R10C25_F5;
assign R10C25_C4 = R10C25_F6;
assign R10C25_C5 = R10C25_F6;
assign R10C25_C6 = R10C25_F4;
assign R10C25_C7 = R10C25_F4;
assign R10C25_N81 = R10C25_Q1;
assign R10C25_S81 = R10C25_Q1;
assign R10C25_E81 = R10C25_Q1;
assign R10C25_W81 = R10C25_Q1;
assign R10C25_N21 = R10C25_Q1;
assign R10C25_N22 = R10C25_Q2;
assign R10C25_S21 = R10C25_Q1;
assign R10C25_S22 = R10C25_Q2;
assign R10C25_E21 = R10C25_Q1;
assign R10C25_E22 = R10C25_Q2;
assign R10C25_W21 = R10C25_Q1;
assign R10C25_W22 = R10C25_Q2;
assign R10C25_E80 = R10C25_Q0;
assign R10C25_W80 = R10C25_Q0;
assign R10C25_N25 = R10C25_Q5;
assign R10C25_N26 = R10C25_Q6;
assign R10C25_S25 = R10C25_Q5;
assign R10C25_S26 = R10C25_Q6;
assign R10C25_N83 = R10C25_Q5;
assign R10C25_S83 = R10C25_Q5;
assign R10C25_N24 = R10C25_Q4;
assign R10C25_N27 = R10C25_Q7;
assign R10C25_S24 = R10C25_Q4;
assign R10C25_S27 = R10C25_Q7;
assign R10C25_N20 = R10C25_Q0;
assign R10C25_N23 = R10C25_Q3;
assign R10C25_S20 = R10C25_Q0;
assign R10C25_S23 = R10C25_Q3;
assign R10C25_N80 = R10C25_Q0;
assign R10C25_S80 = R10C25_Q0;
assign R10C25_E83 = R10C25_Q5;
assign R10C25_W83 = R10C25_Q5;
assign R10C25_E25 = R10C25_Q5;
assign R10C25_E26 = R10C25_Q6;
assign R10C25_W25 = R10C25_Q5;
assign R10C25_W26 = R10C25_Q6;
assign R10C25_E24 = R10C25_Q4;
assign R10C25_E27 = R10C25_Q7;
assign R10C25_W24 = R10C25_Q4;
assign R10C25_W27 = R10C25_Q7;
assign R10C25_E20 = R10C25_Q0;
assign R10C25_E23 = R10C25_Q3;
assign R10C25_W20 = R10C25_Q0;
assign R10C25_W23 = R10C25_Q3;
assign R10C25_B0 = R10C25_F3;
assign R10C25_B1 = R10C25_F3;
assign R10C25_B2 = R10C25_F1;
assign R10C25_B3 = R10C25_F1;
assign R10C25_B4 = R10C25_F1;
assign R10C25_B5 = R10C25_F1;
assign R10C25_B6 = R10C25_F1;
assign R10C25_B7 = R10C25_F1;
assign R10C25_D0 = R10C25_F2;
assign R10C25_D1 = R10C25_F2;
assign R10C25_D2 = R10C25_F0;
assign R10C25_D3 = R10C25_F0;
assign R10C25_D4 = R10C25_F0;
assign R10C25_D5 = R10C25_F0;
assign R10C25_D6 = R10C25_F0;
assign R10C25_D7 = R10C25_F0;
assign R10C25_X02 = R10C25_Q1;
assign R10C25_X04 = R10C25_Q7;
assign R10C25_X06 = R10C25_Q1;
assign R10C25_X08 = R10C25_Q7;
assign R10C25_X01 = R10C25_Q0;
assign R10C25_X03 = R10C25_Q6;
assign R10C25_X05 = R10C25_Q0;
assign R10C25_X07 = R10C25_Q6;
assign R10C25_N10 = R10C25_Q0;
assign R10C25_SN10 = R10C25_Q0;
assign R10C25_SN20 = R10C25_Q0;
assign R10C25_N13 = R10C25_Q0;
assign R10C25_S10 = R10C25_Q0;
assign R10C25_S13 = R10C25_Q0;
assign R10C25_E10 = R10C25_Q0;
assign R10C25_EW10 = R10C25_Q0;
assign R10C25_EW20 = R10C25_Q0;
assign R10C25_E13 = R10C25_Q0;
assign R10C25_W10 = R10C25_Q0;
assign R10C25_W13 = R10C25_Q0;
assign R10C25_E11 = R10C25_EW10;
assign R10C25_W11 = R10C25_EW10;
assign R10C25_E12 = R10C25_EW20;
assign R10C25_W12 = R10C25_EW20;
assign R10C25_S11 = R10C25_SN10;
assign R10C25_N11 = R10C25_SN10;
assign R10C25_S12 = R10C25_SN20;
assign R10C25_N12 = R10C25_SN20;
assign R10C26_CLK0 = VCC;
assign R10C26_CLK1 = VCC;
assign R10C26_CLK2 = VCC;
assign R10C26_LSR0 = VCC;
assign R10C26_LSR1 = VCC;
assign R10C26_LSR2 = VCC;
assign R10C26_CE0 = VCC;
assign R10C26_CE1 = VCC;
assign R10C26_CE2 = VCC;
assign R10C26_SEL0 = VCC;
assign R10C26_SEL1 = VCC;
assign R10C26_SEL2 = VCC;
assign R10C26_SEL3 = VCC;
assign R10C26_SEL4 = VCC;
assign R10C26_SEL5 = VCC;
assign R10C26_SEL6 = VCC;
assign R10C26_SEL7 = VCC;
assign R10C26_C0 = R10C26_F4;
assign R10C26_C1 = R10C26_F4;
assign R10C26_C2 = R10C26_F4;
assign R10C26_C3 = R10C26_F4;
assign R10C26_A4 = R10C26_F7;
assign R10C26_A5 = R10C26_F7;
assign R10C26_A6 = R10C26_F5;
assign R10C26_A7 = R10C26_F5;
assign R10C26_N82 = R10C26_Q4;
assign R10C26_S82 = R10C26_Q4;
assign R10C26_E82 = R10C26_Q4;
assign R10C26_W82 = R10C26_Q4;
assign R10C26_A0 = R10C26_F5;
assign R10C26_A1 = R10C26_F5;
assign R10C26_A2 = R10C26_F5;
assign R10C26_A3 = R10C26_F5;
assign R10C26_C4 = R10C26_F6;
assign R10C26_C5 = R10C26_F6;
assign R10C26_C6 = R10C26_F4;
assign R10C26_C7 = R10C26_F4;
assign R10C26_N81 = R10C26_Q1;
assign R10C26_S81 = R10C26_Q1;
assign R10C26_E81 = R10C26_Q1;
assign R10C26_W81 = R10C26_Q1;
assign R10C26_N21 = R10C26_Q1;
assign R10C26_N22 = R10C26_Q2;
assign R10C26_S21 = R10C26_Q1;
assign R10C26_S22 = R10C26_Q2;
assign R10C26_E21 = R10C26_Q1;
assign R10C26_E22 = R10C26_Q2;
assign R10C26_W21 = R10C26_Q1;
assign R10C26_W22 = R10C26_Q2;
assign R10C26_E80 = R10C26_Q0;
assign R10C26_W80 = R10C26_Q0;
assign R10C26_N25 = R10C26_Q5;
assign R10C26_N26 = R10C26_Q6;
assign R10C26_S25 = R10C26_Q5;
assign R10C26_S26 = R10C26_Q6;
assign R10C26_N83 = R10C26_Q5;
assign R10C26_S83 = R10C26_Q5;
assign R10C26_N24 = R10C26_Q4;
assign R10C26_N27 = R10C26_Q7;
assign R10C26_S24 = R10C26_Q4;
assign R10C26_S27 = R10C26_Q7;
assign R10C26_N20 = R10C26_Q0;
assign R10C26_N23 = R10C26_Q3;
assign R10C26_S20 = R10C26_Q0;
assign R10C26_S23 = R10C26_Q3;
assign R10C26_N80 = R10C26_Q0;
assign R10C26_S80 = R10C26_Q0;
assign R10C26_E83 = R10C26_Q5;
assign R10C26_W83 = R10C26_Q5;
assign R10C26_E25 = R10C26_Q5;
assign R10C26_E26 = R10C26_Q6;
assign R10C26_W25 = R10C26_Q5;
assign R10C26_W26 = R10C26_Q6;
assign R10C26_E24 = R10C26_Q4;
assign R10C26_E27 = R10C26_Q7;
assign R10C26_W24 = R10C26_Q4;
assign R10C26_W27 = R10C26_Q7;
assign R10C26_E20 = R10C26_Q0;
assign R10C26_E23 = R10C26_Q3;
assign R10C26_W20 = R10C26_Q0;
assign R10C26_W23 = R10C26_Q3;
assign R10C26_B0 = R10C26_F3;
assign R10C26_B1 = R10C26_F3;
assign R10C26_B2 = R10C26_F1;
assign R10C26_B3 = R10C26_F1;
assign R10C26_B4 = R10C26_F1;
assign R10C26_B5 = R10C26_F1;
assign R10C26_B6 = R10C26_F1;
assign R10C26_B7 = R10C26_F1;
assign R10C26_D0 = R10C26_F2;
assign R10C26_D1 = R10C26_F2;
assign R10C26_D2 = R10C26_F0;
assign R10C26_D3 = R10C26_F0;
assign R10C26_D4 = R10C26_F0;
assign R10C26_D5 = R10C26_F0;
assign R10C26_D6 = R10C26_F0;
assign R10C26_D7 = R10C26_F0;
assign R10C26_X02 = R10C26_Q1;
assign R10C26_X04 = R10C26_Q7;
assign R10C26_X06 = R10C26_Q1;
assign R10C26_X08 = R10C26_Q7;
assign R10C26_X01 = R10C26_Q0;
assign R10C26_X03 = R10C26_Q6;
assign R10C26_X05 = R10C26_Q0;
assign R10C26_X07 = R10C26_Q6;
assign R10C26_N10 = R10C26_Q0;
assign R10C26_SN10 = R10C26_Q0;
assign R10C26_SN20 = R10C26_Q0;
assign R10C26_N13 = R10C26_Q0;
assign R10C26_S10 = R10C26_Q0;
assign R10C26_S13 = R10C26_Q0;
assign R10C26_E10 = R10C26_Q0;
assign R10C26_EW10 = R10C26_Q0;
assign R10C26_EW20 = R10C26_Q0;
assign R10C26_E13 = R10C26_Q0;
assign R10C26_W10 = R10C26_Q0;
assign R10C26_W13 = R10C26_Q0;
assign R10C26_E11 = R10C26_EW10;
assign R10C26_W11 = R10C26_EW10;
assign R10C26_E12 = R10C26_EW20;
assign R10C26_W12 = R10C26_EW20;
assign R10C26_S11 = R10C26_SN10;
assign R10C26_N11 = R10C26_SN10;
assign R10C26_S12 = R10C26_SN20;
assign R10C26_N12 = R10C26_SN20;
assign R10C27_CLK0 = VCC;
assign R10C27_CLK1 = VCC;
assign R10C27_CLK2 = VCC;
assign R10C27_LSR0 = VCC;
assign R10C27_LSR1 = VCC;
assign R10C27_LSR2 = VCC;
assign R10C27_CE0 = VCC;
assign R10C27_CE1 = VCC;
assign R10C27_CE2 = VCC;
assign R10C27_SEL0 = VCC;
assign R10C27_SEL1 = VCC;
assign R10C27_SEL2 = VCC;
assign R10C27_SEL3 = VCC;
assign R10C27_SEL4 = VCC;
assign R10C27_SEL5 = VCC;
assign R10C27_SEL6 = VCC;
assign R10C27_SEL7 = VCC;
assign R10C27_C0 = R10C27_F4;
assign R10C27_C1 = R10C27_F4;
assign R10C27_C2 = R10C27_F4;
assign R10C27_C3 = R10C27_F4;
assign R10C27_A4 = R10C27_F7;
assign R10C27_A5 = R10C27_F7;
assign R10C27_A6 = R10C27_F5;
assign R10C27_A7 = R10C27_F5;
assign R10C27_N82 = R10C27_Q4;
assign R10C27_S82 = R10C27_Q4;
assign R10C27_E82 = R10C27_Q4;
assign R10C27_W82 = R10C27_Q4;
assign R10C27_A0 = R10C27_F5;
assign R10C27_A1 = R10C27_F5;
assign R10C27_A2 = R10C27_F5;
assign R10C27_A3 = R10C27_F5;
assign R10C27_C4 = R10C27_F6;
assign R10C27_C5 = R10C27_F6;
assign R10C27_C6 = R10C27_F4;
assign R10C27_C7 = R10C27_F4;
assign R10C27_N81 = R10C27_Q1;
assign R10C27_S81 = R10C27_Q1;
assign R10C27_E81 = R10C27_Q1;
assign R10C27_W81 = R10C27_Q1;
assign R10C27_N21 = R10C27_Q1;
assign R10C27_N22 = R10C27_Q2;
assign R10C27_S21 = R10C27_Q1;
assign R10C27_S22 = R10C27_Q2;
assign R10C27_E21 = R10C27_Q1;
assign R10C27_E22 = R10C27_Q2;
assign R10C27_W21 = R10C27_Q1;
assign R10C27_W22 = R10C27_Q2;
assign R10C27_E80 = R10C27_Q0;
assign R10C27_W80 = R10C27_Q0;
assign R10C27_N25 = R10C27_Q5;
assign R10C27_N26 = R10C27_Q6;
assign R10C27_S25 = R10C27_Q5;
assign R10C27_S26 = R10C27_Q6;
assign R10C27_N83 = R10C27_Q5;
assign R10C27_S83 = R10C27_Q5;
assign R10C27_N24 = R10C27_Q4;
assign R10C27_N27 = R10C27_Q7;
assign R10C27_S24 = R10C27_Q4;
assign R10C27_S27 = R10C27_Q7;
assign R10C27_N20 = R10C27_Q0;
assign R10C27_N23 = R10C27_Q3;
assign R10C27_S20 = R10C27_Q0;
assign R10C27_S23 = R10C27_Q3;
assign R10C27_N80 = R10C27_Q0;
assign R10C27_S80 = R10C27_Q0;
assign R10C27_E83 = R10C27_Q5;
assign R10C27_W83 = R10C27_Q5;
assign R10C27_E25 = R10C27_Q5;
assign R10C27_E26 = R10C27_Q6;
assign R10C27_W25 = R10C27_Q5;
assign R10C27_W26 = R10C27_Q6;
assign R10C27_E24 = R10C27_Q4;
assign R10C27_E27 = R10C27_Q7;
assign R10C27_W24 = R10C27_Q4;
assign R10C27_W27 = R10C27_Q7;
assign R10C27_E20 = R10C27_Q0;
assign R10C27_E23 = R10C27_Q3;
assign R10C27_W20 = R10C27_Q0;
assign R10C27_W23 = R10C27_Q3;
assign R10C27_B0 = R10C27_F3;
assign R10C27_B1 = R10C27_F3;
assign R10C27_B2 = R10C27_F1;
assign R10C27_B3 = R10C27_F1;
assign R10C27_B4 = R10C27_F1;
assign R10C27_B5 = R10C27_F1;
assign R10C27_B6 = R10C27_F1;
assign R10C27_B7 = R10C27_F1;
assign R10C27_D0 = R10C27_F2;
assign R10C27_D1 = R10C27_F2;
assign R10C27_D2 = R10C27_F0;
assign R10C27_D3 = R10C27_F0;
assign R10C27_D4 = R10C27_F0;
assign R10C27_D5 = R10C27_F0;
assign R10C27_D6 = R10C27_F0;
assign R10C27_D7 = R10C27_F0;
assign R10C27_X02 = R10C27_Q1;
assign R10C27_X04 = R10C27_Q7;
assign R10C27_X06 = R10C27_Q1;
assign R10C27_X08 = R10C27_Q7;
assign R10C27_X01 = R10C27_Q0;
assign R10C27_X03 = R10C27_Q6;
assign R10C27_X05 = R10C27_Q0;
assign R10C27_X07 = R10C27_Q6;
assign R10C27_N10 = R10C27_Q0;
assign R10C27_SN10 = R10C27_Q0;
assign R10C27_SN20 = R10C27_Q0;
assign R10C27_N13 = R10C27_Q0;
assign R10C27_S10 = R10C27_Q0;
assign R10C27_S13 = R10C27_Q0;
assign R10C27_E10 = R10C27_Q0;
assign R10C27_EW10 = R10C27_Q0;
assign R10C27_EW20 = R10C27_Q0;
assign R10C27_E13 = R10C27_Q0;
assign R10C27_W10 = R10C27_Q0;
assign R10C27_W13 = R10C27_Q0;
assign R10C27_E11 = R10C27_EW10;
assign R10C27_W11 = R10C27_EW10;
assign R10C27_E12 = R10C27_EW20;
assign R10C27_W12 = R10C27_EW20;
assign R10C27_S11 = R10C27_SN10;
assign R10C27_N11 = R10C27_SN10;
assign R10C27_S12 = R10C27_SN20;
assign R10C27_N12 = R10C27_SN20;
assign R10C28_CLK0 = VCC;
assign R10C28_CLK1 = VCC;
assign R10C28_CLK2 = VCC;
assign R10C28_LSR0 = VCC;
assign R10C28_LSR1 = VCC;
assign R10C28_LSR2 = VCC;
assign R10C28_CE0 = VCC;
assign R10C28_CE1 = VCC;
assign R10C28_CE2 = VCC;
assign R10C28_SEL0 = VCC;
assign R10C28_SEL1 = VCC;
assign R10C28_SEL2 = VCC;
assign R10C28_SEL3 = VCC;
assign R10C28_SEL4 = VCC;
assign R10C28_SEL5 = VCC;
assign R10C28_SEL6 = VCC;
assign R10C28_SEL7 = VCC;
assign R10C28_C0 = R10C28_F4;
assign R10C28_C1 = R10C28_F4;
assign R10C28_C2 = R10C28_F4;
assign R10C28_C3 = R10C28_F4;
assign R10C28_A4 = R10C28_F7;
assign R10C28_A5 = R10C28_F7;
assign R10C28_A6 = R10C28_F5;
assign R10C28_A7 = R10C28_F5;
assign R10C28_N82 = R10C28_Q4;
assign R10C28_S82 = R10C28_Q4;
assign R10C28_E82 = R10C28_Q4;
assign R10C28_W82 = R10C28_Q4;
assign R10C28_A0 = R10C28_F5;
assign R10C28_A1 = R10C28_F5;
assign R10C28_A2 = R10C28_F5;
assign R10C28_A3 = R10C28_F5;
assign R10C28_C4 = R10C28_F6;
assign R10C28_C5 = R10C28_F6;
assign R10C28_C6 = R10C28_F4;
assign R10C28_C7 = R10C28_F4;
assign R10C28_N81 = R10C28_Q1;
assign R10C28_S81 = R10C28_Q1;
assign R10C28_E81 = R10C28_Q1;
assign R10C28_W81 = R10C28_Q1;
assign R10C28_N21 = R10C28_Q1;
assign R10C28_N22 = R10C28_Q2;
assign R10C28_S21 = R10C28_Q1;
assign R10C28_S22 = R10C28_Q2;
assign R10C28_E21 = R10C28_Q1;
assign R10C28_E22 = R10C28_Q2;
assign R10C28_W21 = R10C28_Q1;
assign R10C28_W22 = R10C28_Q2;
assign R10C28_E80 = R10C28_Q0;
assign R10C28_W80 = R10C28_Q0;
assign R10C28_N25 = R10C28_Q5;
assign R10C28_N26 = R10C28_Q6;
assign R10C28_S25 = R10C28_Q5;
assign R10C28_S26 = R10C28_Q6;
assign R10C28_N83 = R10C28_Q5;
assign R10C28_S83 = R10C28_Q5;
assign R10C28_N24 = R10C28_Q4;
assign R10C28_N27 = R10C28_Q7;
assign R10C28_S24 = R10C28_Q4;
assign R10C28_S27 = R10C28_Q7;
assign R10C28_N20 = R10C28_Q0;
assign R10C28_N23 = R10C28_Q3;
assign R10C28_S20 = R10C28_Q0;
assign R10C28_S23 = R10C28_Q3;
assign R10C28_N80 = R10C28_Q0;
assign R10C28_S80 = R10C28_Q0;
assign R10C28_E83 = R10C28_Q5;
assign R10C28_W83 = R10C28_Q5;
assign R10C28_E25 = R10C28_Q5;
assign R10C28_E26 = R10C28_Q6;
assign R10C28_W25 = R10C28_Q5;
assign R10C28_W26 = R10C28_Q6;
assign R10C28_E24 = R10C28_Q4;
assign R10C28_E27 = R10C28_Q7;
assign R10C28_W24 = R10C28_Q4;
assign R10C28_W27 = R10C28_Q7;
assign R10C28_E20 = R10C28_Q0;
assign R10C28_E23 = R10C28_Q3;
assign R10C28_W20 = R10C28_Q0;
assign R10C28_W23 = R10C28_Q3;
assign R10C28_B0 = R10C28_F3;
assign R10C28_B1 = R10C28_F3;
assign R10C28_B2 = R10C28_F1;
assign R10C28_B3 = R10C28_F1;
assign R10C28_B4 = R10C28_F1;
assign R10C28_B5 = R10C28_F1;
assign R10C28_B6 = R10C28_F1;
assign R10C28_B7 = R10C28_F1;
assign R10C28_D0 = R10C28_F2;
assign R10C28_D1 = R10C28_F2;
assign R10C28_D2 = R10C28_F0;
assign R10C28_D3 = R10C28_F0;
assign R10C28_D4 = R10C28_F0;
assign R10C28_D5 = R10C28_F0;
assign R10C28_D6 = R10C28_F0;
assign R10C28_D7 = R10C28_F0;
assign R10C28_X02 = R10C28_Q1;
assign R10C28_X04 = R10C28_Q7;
assign R10C28_X06 = R10C28_Q1;
assign R10C28_X08 = R10C28_Q7;
assign R10C28_X01 = R10C28_Q0;
assign R10C28_X03 = R10C28_Q6;
assign R10C28_X05 = R10C28_Q0;
assign R10C28_X07 = R10C28_Q6;
assign R10C28_N10 = R10C28_Q0;
assign R10C28_SN10 = R10C28_Q0;
assign R10C28_SN20 = R10C28_Q0;
assign R10C28_N13 = R10C28_Q0;
assign R10C28_S10 = R10C28_Q0;
assign R10C28_S13 = R10C28_Q0;
assign R10C28_E10 = R10C28_Q0;
assign R10C28_EW10 = R10C28_Q0;
assign R10C28_EW20 = R10C28_Q0;
assign R10C28_E13 = R10C28_Q0;
assign R10C28_W10 = R10C28_Q0;
assign R10C28_W13 = R10C28_Q0;
assign R10C28_E11 = R10C28_EW10;
assign R10C28_W11 = R10C28_EW10;
assign R10C28_E12 = R10C28_EW20;
assign R10C28_W12 = R10C28_EW20;
assign R10C28_S11 = R10C28_SN10;
assign R10C28_N11 = R10C28_SN10;
assign R10C28_S12 = R10C28_SN20;
assign R10C28_N12 = R10C28_SN20;
assign R10C29_CLK0 = VCC;
assign R10C29_CLK1 = VCC;
assign R10C29_CLK2 = VCC;
assign R10C29_LSR0 = VCC;
assign R10C29_LSR1 = VCC;
assign R10C29_LSR2 = VCC;
assign R10C29_CE0 = VCC;
assign R10C29_CE1 = VCC;
assign R10C29_CE2 = VCC;
assign R10C29_SEL0 = VCC;
assign R10C29_SEL1 = VCC;
assign R10C29_SEL2 = VCC;
assign R10C29_SEL3 = VCC;
assign R10C29_SEL4 = VCC;
assign R10C29_SEL5 = VCC;
assign R10C29_SEL6 = VCC;
assign R10C29_SEL7 = VCC;
assign R10C29_C0 = R10C29_F4;
assign R10C29_C1 = R10C29_F4;
assign R10C29_C2 = R10C29_F4;
assign R10C29_C3 = R10C29_F4;
assign R10C29_A4 = R10C29_F7;
assign R10C29_A5 = R10C29_F7;
assign R10C29_A6 = R10C29_F5;
assign R10C29_A7 = R10C29_F5;
assign R10C29_N82 = R10C29_Q4;
assign R10C29_S82 = R10C29_Q4;
assign R10C29_E82 = R10C29_Q4;
assign R10C29_W82 = R10C29_Q4;
assign R10C29_A0 = R10C29_F5;
assign R10C29_A1 = R10C29_F5;
assign R10C29_A2 = R10C29_F5;
assign R10C29_A3 = R10C29_F5;
assign R10C29_C4 = R10C29_F6;
assign R10C29_C5 = R10C29_F6;
assign R10C29_C6 = R10C29_F4;
assign R10C29_C7 = R10C29_F4;
assign R10C29_N81 = R10C29_Q1;
assign R10C29_S81 = R10C29_Q1;
assign R10C29_E81 = R10C29_Q1;
assign R10C29_W81 = R10C29_Q1;
assign R10C29_N21 = R10C29_Q1;
assign R10C29_N22 = R10C29_Q2;
assign R10C29_S21 = R10C29_Q1;
assign R10C29_S22 = R10C29_Q2;
assign R10C29_E21 = R10C29_Q1;
assign R10C29_E22 = R10C29_Q2;
assign R10C29_W21 = R10C29_Q1;
assign R10C29_W22 = R10C29_Q2;
assign R10C29_E80 = R10C29_Q0;
assign R10C29_W80 = R10C29_Q0;
assign R10C29_N25 = R10C29_Q5;
assign R10C29_N26 = R10C29_Q6;
assign R10C29_S25 = R10C29_Q5;
assign R10C29_S26 = R10C29_Q6;
assign R10C29_N83 = R10C29_Q5;
assign R10C29_S83 = R10C29_Q5;
assign R10C29_N24 = R10C29_Q4;
assign R10C29_N27 = R10C29_Q7;
assign R10C29_S24 = R10C29_Q4;
assign R10C29_S27 = R10C29_Q7;
assign R10C29_N20 = R10C29_Q0;
assign R10C29_N23 = R10C29_Q3;
assign R10C29_S20 = R10C29_Q0;
assign R10C29_S23 = R10C29_Q3;
assign R10C29_N80 = R10C29_Q0;
assign R10C29_S80 = R10C29_Q0;
assign R10C29_E83 = R10C29_Q5;
assign R10C29_W83 = R10C29_Q5;
assign R10C29_E25 = R10C29_Q5;
assign R10C29_E26 = R10C29_Q6;
assign R10C29_W25 = R10C29_Q5;
assign R10C29_W26 = R10C29_Q6;
assign R10C29_E24 = R10C29_Q4;
assign R10C29_E27 = R10C29_Q7;
assign R10C29_W24 = R10C29_Q4;
assign R10C29_W27 = R10C29_Q7;
assign R10C29_E20 = R10C29_Q0;
assign R10C29_E23 = R10C29_Q3;
assign R10C29_W20 = R10C29_Q0;
assign R10C29_W23 = R10C29_Q3;
assign R10C29_B0 = R10C29_F3;
assign R10C29_B1 = R10C29_F3;
assign R10C29_B2 = R10C29_F1;
assign R10C29_B3 = R10C29_F1;
assign R10C29_B4 = R10C29_F1;
assign R10C29_B5 = R10C29_F1;
assign R10C29_B6 = R10C29_F1;
assign R10C29_B7 = R10C29_F1;
assign R10C29_D0 = R10C29_F2;
assign R10C29_D1 = R10C29_F2;
assign R10C29_D2 = R10C29_F0;
assign R10C29_D3 = R10C29_F0;
assign R10C29_D4 = R10C29_F0;
assign R10C29_D5 = R10C29_F0;
assign R10C29_D6 = R10C29_F0;
assign R10C29_D7 = R10C29_F0;
assign R10C29_X02 = R10C29_Q1;
assign R10C29_X04 = R10C29_Q7;
assign R10C29_X06 = R10C29_Q1;
assign R10C29_X08 = R10C29_Q7;
assign R10C29_X01 = R10C29_Q0;
assign R10C29_X03 = R10C29_Q6;
assign R10C29_X05 = R10C29_Q0;
assign R10C29_X07 = R10C29_Q6;
assign R10C29_N10 = R10C29_Q0;
assign R10C29_SN10 = R10C29_Q0;
assign R10C29_SN20 = R10C29_Q0;
assign R10C29_N13 = R10C29_Q0;
assign R10C29_S10 = R10C29_Q0;
assign R10C29_S13 = R10C29_Q0;
assign R10C29_E10 = R10C29_Q0;
assign R10C29_EW10 = R10C29_Q0;
assign R10C29_EW20 = R10C29_Q0;
assign R10C29_E13 = R10C29_Q0;
assign R10C29_W10 = R10C29_Q0;
assign R10C29_W13 = R10C29_Q0;
assign R10C29_E11 = R10C29_EW10;
assign R10C29_W11 = R10C29_EW10;
assign R10C29_E12 = R10C29_EW20;
assign R10C29_W12 = R10C29_EW20;
assign R10C29_S11 = R10C29_SN10;
assign R10C29_N11 = R10C29_SN10;
assign R10C29_S12 = R10C29_SN20;
assign R10C29_N12 = R10C29_SN20;
assign R10C30_CLK0 = VCC;
assign R10C30_CLK1 = VCC;
assign R10C30_CLK2 = VCC;
assign R10C30_LSR0 = VCC;
assign R10C30_LSR1 = VCC;
assign R10C30_LSR2 = VCC;
assign R10C30_CE0 = VCC;
assign R10C30_CE1 = VCC;
assign R10C30_CE2 = VCC;
assign R10C30_SEL0 = VCC;
assign R10C30_SEL1 = VCC;
assign R10C30_SEL2 = VCC;
assign R10C30_SEL3 = VCC;
assign R10C30_SEL4 = VCC;
assign R10C30_SEL5 = VCC;
assign R10C30_SEL6 = VCC;
assign R10C30_SEL7 = VCC;
assign R10C30_C0 = R10C30_F4;
assign R10C30_C1 = R10C30_F4;
assign R10C30_C2 = R10C30_F4;
assign R10C30_C3 = R10C30_F4;
assign R10C30_A4 = R10C30_F7;
assign R10C30_A5 = R10C30_F7;
assign R10C30_A6 = R10C30_F5;
assign R10C30_A7 = R10C30_F5;
assign R10C30_N82 = R10C30_Q4;
assign R10C30_S82 = R10C30_Q4;
assign R10C30_E82 = R10C30_Q4;
assign R10C30_W82 = R10C30_Q4;
assign R10C30_A0 = R10C30_F5;
assign R10C30_A1 = R10C30_F5;
assign R10C30_A2 = R10C30_F5;
assign R10C30_A3 = R10C30_F5;
assign R10C30_C4 = R10C30_F6;
assign R10C30_C5 = R10C30_F6;
assign R10C30_C6 = R10C30_F4;
assign R10C30_C7 = R10C30_F4;
assign R10C30_N81 = R10C30_Q1;
assign R10C30_S81 = R10C30_Q1;
assign R10C30_E81 = R10C30_Q1;
assign R10C30_W81 = R10C30_Q1;
assign R10C30_N21 = R10C30_Q1;
assign R10C30_N22 = R10C30_Q2;
assign R10C30_S21 = R10C30_Q1;
assign R10C30_S22 = R10C30_Q2;
assign R10C30_E21 = R10C30_Q1;
assign R10C30_E22 = R10C30_Q2;
assign R10C30_W21 = R10C30_Q1;
assign R10C30_W22 = R10C30_Q2;
assign R10C30_E80 = R10C30_Q0;
assign R10C30_W80 = R10C30_Q0;
assign R10C30_N25 = R10C30_Q5;
assign R10C30_N26 = R10C30_Q6;
assign R10C30_S25 = R10C30_Q5;
assign R10C30_S26 = R10C30_Q6;
assign R10C30_N83 = R10C30_Q5;
assign R10C30_S83 = R10C30_Q5;
assign R10C30_N24 = R10C30_Q4;
assign R10C30_N27 = R10C30_Q7;
assign R10C30_S24 = R10C30_Q4;
assign R10C30_S27 = R10C30_Q7;
assign R10C30_N20 = R10C30_Q0;
assign R10C30_N23 = R10C30_Q3;
assign R10C30_S20 = R10C30_Q0;
assign R10C30_S23 = R10C30_Q3;
assign R10C30_N80 = R10C30_Q0;
assign R10C30_S80 = R10C30_Q0;
assign R10C30_E83 = R10C30_Q5;
assign R10C30_W83 = R10C30_Q5;
assign R10C30_E25 = R10C30_Q5;
assign R10C30_E26 = R10C30_Q6;
assign R10C30_W25 = R10C30_Q5;
assign R10C30_W26 = R10C30_Q6;
assign R10C30_E24 = R10C30_Q4;
assign R10C30_E27 = R10C30_Q7;
assign R10C30_W24 = R10C30_Q4;
assign R10C30_W27 = R10C30_Q7;
assign R10C30_E20 = R10C30_Q0;
assign R10C30_E23 = R10C30_Q3;
assign R10C30_W20 = R10C30_Q0;
assign R10C30_W23 = R10C30_Q3;
assign R10C30_B0 = R10C30_F3;
assign R10C30_B1 = R10C30_F3;
assign R10C30_B2 = R10C30_F1;
assign R10C30_B3 = R10C30_F1;
assign R10C30_B4 = R10C30_F1;
assign R10C30_B5 = R10C30_F1;
assign R10C30_B6 = R10C30_F1;
assign R10C30_B7 = R10C30_F1;
assign R10C30_D0 = R10C30_F2;
assign R10C30_D1 = R10C30_F2;
assign R10C30_D2 = R10C30_F0;
assign R10C30_D3 = R10C30_F0;
assign R10C30_D4 = R10C30_F0;
assign R10C30_D5 = R10C30_F0;
assign R10C30_D6 = R10C30_F0;
assign R10C30_D7 = R10C30_F0;
assign R10C30_X02 = R10C30_Q1;
assign R10C30_X04 = R10C30_Q7;
assign R10C30_X06 = R10C30_Q1;
assign R10C30_X08 = R10C30_Q7;
assign R10C30_X01 = R10C30_Q0;
assign R10C30_X03 = R10C30_Q6;
assign R10C30_X05 = R10C30_Q0;
assign R10C30_X07 = R10C30_Q6;
assign R10C30_N10 = R10C30_Q0;
assign R10C30_SN10 = R10C30_Q0;
assign R10C30_SN20 = R10C30_Q0;
assign R10C30_N13 = R10C30_Q0;
assign R10C30_S10 = R10C30_Q0;
assign R10C30_S13 = R10C30_Q0;
assign R10C30_E10 = R10C30_Q0;
assign R10C30_EW10 = R10C30_Q0;
assign R10C30_EW20 = R10C30_Q0;
assign R10C30_E13 = R10C30_Q0;
assign R10C30_W10 = R10C30_Q0;
assign R10C30_W13 = R10C30_Q0;
assign R10C30_E11 = R10C30_EW10;
assign R10C30_W11 = R10C30_EW10;
assign R10C30_E12 = R10C30_EW20;
assign R10C30_W12 = R10C30_EW20;
assign R10C30_S11 = R10C30_SN10;
assign R10C30_N11 = R10C30_SN10;
assign R10C30_S12 = R10C30_SN20;
assign R10C30_N12 = R10C30_SN20;
assign R10C31_CLK0 = VCC;
assign R10C31_CLK1 = VCC;
assign R10C31_CLK2 = VCC;
assign R10C31_LSR0 = VCC;
assign R10C31_LSR1 = VCC;
assign R10C31_LSR2 = VCC;
assign R10C31_CE0 = VCC;
assign R10C31_CE1 = VCC;
assign R10C31_CE2 = VCC;
assign R10C31_SEL0 = VCC;
assign R10C31_SEL1 = VCC;
assign R10C31_SEL2 = VCC;
assign R10C31_SEL3 = VCC;
assign R10C31_SEL4 = VCC;
assign R10C31_SEL5 = VCC;
assign R10C31_SEL6 = VCC;
assign R10C31_SEL7 = VCC;
assign R10C31_C0 = R10C31_F4;
assign R10C31_C1 = R10C31_F4;
assign R10C31_C2 = R10C31_F4;
assign R10C31_C3 = R10C31_F4;
assign R10C31_A4 = R10C31_F7;
assign R10C31_A5 = R10C31_F7;
assign R10C31_A6 = R10C31_F5;
assign R10C31_A7 = R10C31_F5;
assign R10C31_N82 = R10C31_Q4;
assign R10C31_S82 = R10C31_Q4;
assign R10C31_E82 = R10C31_Q4;
assign R10C31_W82 = R10C31_Q4;
assign R10C31_A0 = R10C31_F5;
assign R10C31_A1 = R10C31_F5;
assign R10C31_A2 = R10C31_F5;
assign R10C31_A3 = R10C31_F5;
assign R10C31_C4 = R10C31_F6;
assign R10C31_C5 = R10C31_F6;
assign R10C31_C6 = R10C31_F4;
assign R10C31_C7 = R10C31_F4;
assign R10C31_N81 = R10C31_Q1;
assign R10C31_S81 = R10C31_Q1;
assign R10C31_E81 = R10C31_Q1;
assign R10C31_W81 = R10C31_Q1;
assign R10C31_N21 = R10C31_Q1;
assign R10C31_N22 = R10C31_Q2;
assign R10C31_S21 = R10C31_Q1;
assign R10C31_S22 = R10C31_Q2;
assign R10C31_E21 = R10C31_Q1;
assign R10C31_E22 = R10C31_Q2;
assign R10C31_W21 = R10C31_Q1;
assign R10C31_W22 = R10C31_Q2;
assign R10C31_E80 = R10C31_Q0;
assign R10C31_W80 = R10C31_Q0;
assign R10C31_N25 = R10C31_Q5;
assign R10C31_N26 = R10C31_Q6;
assign R10C31_S25 = R10C31_Q5;
assign R10C31_S26 = R10C31_Q6;
assign R10C31_N83 = R10C31_Q5;
assign R10C31_S83 = R10C31_Q5;
assign R10C31_N24 = R10C31_Q4;
assign R10C31_N27 = R10C31_Q7;
assign R10C31_S24 = R10C31_Q4;
assign R10C31_S27 = R10C31_Q7;
assign R10C31_N20 = R10C31_Q0;
assign R10C31_N23 = R10C31_Q3;
assign R10C31_S20 = R10C31_Q0;
assign R10C31_S23 = R10C31_Q3;
assign R10C31_N80 = R10C31_Q0;
assign R10C31_S80 = R10C31_Q0;
assign R10C31_E83 = R10C31_Q5;
assign R10C31_W83 = R10C31_Q5;
assign R10C31_E25 = R10C31_Q5;
assign R10C31_E26 = R10C31_Q6;
assign R10C31_W25 = R10C31_Q5;
assign R10C31_W26 = R10C31_Q6;
assign R10C31_E24 = R10C31_Q4;
assign R10C31_E27 = R10C31_Q7;
assign R10C31_W24 = R10C31_Q4;
assign R10C31_W27 = R10C31_Q7;
assign R10C31_E20 = R10C31_Q0;
assign R10C31_E23 = R10C31_Q3;
assign R10C31_W20 = R10C31_Q0;
assign R10C31_W23 = R10C31_Q3;
assign R10C31_B0 = R10C31_F3;
assign R10C31_B1 = R10C31_F3;
assign R10C31_B2 = R10C31_F1;
assign R10C31_B3 = R10C31_F1;
assign R10C31_B4 = R10C31_F1;
assign R10C31_B5 = R10C31_F1;
assign R10C31_B6 = R10C31_F1;
assign R10C31_B7 = R10C31_F1;
assign R10C31_D0 = R10C31_F2;
assign R10C31_D1 = R10C31_F2;
assign R10C31_D2 = R10C31_F0;
assign R10C31_D3 = R10C31_F0;
assign R10C31_D4 = R10C31_F0;
assign R10C31_D5 = R10C31_F0;
assign R10C31_D6 = R10C31_F0;
assign R10C31_D7 = R10C31_F0;
assign R10C31_X02 = R10C31_Q1;
assign R10C31_X04 = R10C31_Q7;
assign R10C31_X06 = R10C31_Q1;
assign R10C31_X08 = R10C31_Q7;
assign R10C31_X01 = R10C31_Q0;
assign R10C31_X03 = R10C31_Q6;
assign R10C31_X05 = R10C31_Q0;
assign R10C31_X07 = R10C31_Q6;
assign R10C31_N10 = R10C31_Q0;
assign R10C31_SN10 = R10C31_Q0;
assign R10C31_SN20 = R10C31_Q0;
assign R10C31_N13 = R10C31_Q0;
assign R10C31_S10 = R10C31_Q0;
assign R10C31_S13 = R10C31_Q0;
assign R10C31_E10 = R10C31_Q0;
assign R10C31_EW10 = R10C31_Q0;
assign R10C31_EW20 = R10C31_Q0;
assign R10C31_E13 = R10C31_Q0;
assign R10C31_W10 = R10C31_Q0;
assign R10C31_W13 = R10C31_Q0;
assign R10C31_E11 = R10C31_EW10;
assign R10C31_W11 = R10C31_EW10;
assign R10C31_E12 = R10C31_EW20;
assign R10C31_W12 = R10C31_EW20;
assign R10C31_S11 = R10C31_SN10;
assign R10C31_N11 = R10C31_SN10;
assign R10C31_S12 = R10C31_SN20;
assign R10C31_N12 = R10C31_SN20;
assign R10C34_CLK0 = VCC;
assign R10C34_CLK1 = VCC;
assign R10C34_CLK2 = VCC;
assign R10C34_LSR0 = VCC;
assign R10C34_LSR1 = VCC;
assign R10C34_LSR2 = VCC;
assign R10C34_CE0 = VCC;
assign R10C34_CE1 = VCC;
assign R10C34_CE2 = VCC;
assign R10C34_SEL0 = VCC;
assign R10C34_SEL1 = VCC;
assign R10C34_SEL2 = VCC;
assign R10C34_SEL3 = VCC;
assign R10C34_SEL4 = VCC;
assign R10C34_SEL5 = VCC;
assign R10C34_SEL6 = VCC;
assign R10C34_SEL7 = VCC;
assign R10C34_C0 = R10C34_F4;
assign R10C34_C1 = R10C34_F4;
assign R10C34_C2 = R10C34_F4;
assign R10C34_C3 = R10C34_F4;
assign R10C34_A4 = R10C34_F7;
assign R10C34_A5 = R10C34_F7;
assign R10C34_A6 = R10C34_F5;
assign R10C34_A7 = R10C34_F5;
assign R10C34_N82 = R10C34_Q4;
assign R10C34_S82 = R10C34_Q4;
assign R10C34_E82 = R10C34_Q4;
assign R10C34_W82 = R10C34_Q4;
assign R10C34_A0 = R10C34_F5;
assign R10C34_A1 = R10C34_F5;
assign R10C34_A2 = R10C34_F5;
assign R10C34_A3 = R10C34_F5;
assign R10C34_C4 = R10C34_F6;
assign R10C34_C5 = R10C34_F6;
assign R10C34_C6 = R10C34_F4;
assign R10C34_C7 = R10C34_F4;
assign R10C34_N81 = R10C34_Q1;
assign R10C34_S81 = R10C34_Q1;
assign R10C34_E81 = R10C34_Q1;
assign R10C34_W81 = R10C34_Q1;
assign R10C34_N21 = R10C34_Q1;
assign R10C34_N22 = R10C34_Q2;
assign R10C34_S21 = R10C34_Q1;
assign R10C34_S22 = R10C34_Q2;
assign R10C34_E21 = R10C34_Q1;
assign R10C34_E22 = R10C34_Q2;
assign R10C34_W21 = R10C34_Q1;
assign R10C34_W22 = R10C34_Q2;
assign R10C34_E80 = R10C34_Q0;
assign R10C34_W80 = R10C34_Q0;
assign R10C34_N25 = R10C34_Q5;
assign R10C34_N26 = R10C34_Q6;
assign R10C34_S25 = R10C34_Q5;
assign R10C34_S26 = R10C34_Q6;
assign R10C34_N83 = R10C34_Q5;
assign R10C34_S83 = R10C34_Q5;
assign R10C34_N24 = R10C34_Q4;
assign R10C34_N27 = R10C34_Q7;
assign R10C34_S24 = R10C34_Q4;
assign R10C34_S27 = R10C34_Q7;
assign R10C34_N20 = R10C34_Q0;
assign R10C34_N23 = R10C34_Q3;
assign R10C34_S20 = R10C34_Q0;
assign R10C34_S23 = R10C34_Q3;
assign R10C34_N80 = R10C34_Q0;
assign R10C34_S80 = R10C34_Q0;
assign R10C34_E83 = R10C34_Q5;
assign R10C34_W83 = R10C34_Q5;
assign R10C34_E25 = R10C34_Q5;
assign R10C34_E26 = R10C34_Q6;
assign R10C34_W25 = R10C34_Q5;
assign R10C34_W26 = R10C34_Q6;
assign R10C34_E24 = R10C34_Q4;
assign R10C34_E27 = R10C34_Q7;
assign R10C34_W24 = R10C34_Q4;
assign R10C34_W27 = R10C34_Q7;
assign R10C34_E20 = R10C34_Q0;
assign R10C34_E23 = R10C34_Q3;
assign R10C34_W20 = R10C34_Q0;
assign R10C34_W23 = R10C34_Q3;
assign R10C34_B0 = R10C34_F3;
assign R10C34_B1 = R10C34_F3;
assign R10C34_B2 = R10C34_F1;
assign R10C34_B3 = R10C34_F1;
assign R10C34_B4 = R10C34_F1;
assign R10C34_B5 = R10C34_F1;
assign R10C34_B6 = R10C34_F1;
assign R10C34_B7 = R10C34_F1;
assign R10C34_D0 = R10C34_F2;
assign R10C34_D1 = R10C34_F2;
assign R10C34_D2 = R10C34_F0;
assign R10C34_D3 = R10C34_F0;
assign R10C34_D4 = R10C34_F0;
assign R10C34_D5 = R10C34_F0;
assign R10C34_D6 = R10C34_F0;
assign R10C34_D7 = R10C34_F0;
assign R10C34_X02 = R10C34_Q1;
assign R10C34_X04 = R10C34_Q7;
assign R10C34_X06 = R10C34_Q1;
assign R10C34_X08 = R10C34_Q7;
assign R10C34_X01 = R10C34_Q0;
assign R10C34_X03 = R10C34_Q6;
assign R10C34_X05 = R10C34_Q0;
assign R10C34_X07 = R10C34_Q6;
assign R10C34_N10 = R10C34_Q0;
assign R10C34_SN10 = R10C34_Q0;
assign R10C34_SN20 = R10C34_Q0;
assign R10C34_N13 = R10C34_Q0;
assign R10C34_S10 = R10C34_Q0;
assign R10C34_S13 = R10C34_Q0;
assign R10C34_E10 = R10C34_Q0;
assign R10C34_EW10 = R10C34_Q0;
assign R10C34_EW20 = R10C34_Q0;
assign R10C34_E13 = R10C34_Q0;
assign R10C34_W10 = R10C34_Q0;
assign R10C34_W13 = R10C34_Q0;
assign R10C34_E11 = R10C34_EW10;
assign R10C34_W11 = R10C34_EW10;
assign R10C34_E12 = R10C34_EW20;
assign R10C34_W12 = R10C34_EW20;
assign R10C34_S11 = R10C34_SN10;
assign R10C34_N11 = R10C34_SN10;
assign R10C34_S12 = R10C34_SN20;
assign R10C34_N12 = R10C34_SN20;
assign R10C37_CLK0 = VCC;
assign R10C37_CLK1 = VCC;
assign R10C37_CLK2 = VCC;
assign R10C37_LSR0 = VCC;
assign R10C37_LSR1 = VCC;
assign R10C37_LSR2 = VCC;
assign R10C37_CE0 = VCC;
assign R10C37_CE1 = VCC;
assign R10C37_CE2 = VCC;
assign R10C37_SEL0 = VCC;
assign R10C37_SEL1 = VCC;
assign R10C37_SEL2 = VCC;
assign R10C37_SEL3 = VCC;
assign R10C37_SEL4 = VCC;
assign R10C37_SEL5 = VCC;
assign R10C37_SEL6 = VCC;
assign R10C37_SEL7 = VCC;
assign R10C37_C0 = R10C37_F4;
assign R10C37_C1 = R10C37_F4;
assign R10C37_C2 = R10C37_F4;
assign R10C37_C3 = R10C37_F4;
assign R10C37_A4 = R10C37_F7;
assign R10C37_A5 = R10C37_F7;
assign R10C37_A6 = R10C37_F5;
assign R10C37_A7 = R10C37_F5;
assign R10C37_N82 = R10C37_Q4;
assign R10C37_S82 = R10C37_Q4;
assign R10C37_E82 = R10C37_Q4;
assign R10C37_W82 = R10C37_Q4;
assign R10C37_A0 = R10C37_F5;
assign R10C37_A1 = R10C37_F5;
assign R10C37_A2 = R10C37_F5;
assign R10C37_A3 = R10C37_F5;
assign R10C37_C4 = R10C37_F6;
assign R10C37_C5 = R10C37_F6;
assign R10C37_C6 = R10C37_F4;
assign R10C37_C7 = R10C37_F4;
assign R10C37_N81 = R10C37_Q1;
assign R10C37_S81 = R10C37_Q1;
assign R10C37_E81 = R10C37_Q1;
assign R10C37_W81 = R10C37_Q1;
assign R10C37_N21 = R10C37_Q1;
assign R10C37_N22 = R10C37_Q2;
assign R10C37_S21 = R10C37_Q1;
assign R10C37_S22 = R10C37_Q2;
assign R10C37_E21 = R10C37_Q1;
assign R10C37_E22 = R10C37_Q2;
assign R10C37_W21 = R10C37_Q1;
assign R10C37_W22 = R10C37_Q2;
assign R10C37_E80 = R10C37_Q0;
assign R10C37_W80 = R10C37_Q0;
assign R10C37_N25 = R10C37_Q5;
assign R10C37_N26 = R10C37_Q6;
assign R10C37_S25 = R10C37_Q5;
assign R10C37_S26 = R10C37_Q6;
assign R10C37_N83 = R10C37_Q5;
assign R10C37_S83 = R10C37_Q5;
assign R10C37_N24 = R10C37_Q4;
assign R10C37_N27 = R10C37_Q7;
assign R10C37_S24 = R10C37_Q4;
assign R10C37_S27 = R10C37_Q7;
assign R10C37_N20 = R10C37_Q0;
assign R10C37_N23 = R10C37_Q3;
assign R10C37_S20 = R10C37_Q0;
assign R10C37_S23 = R10C37_Q3;
assign R10C37_N80 = R10C37_Q0;
assign R10C37_S80 = R10C37_Q0;
assign R10C37_E83 = R10C37_Q5;
assign R10C37_W83 = R10C37_Q5;
assign R10C37_E25 = R10C37_Q5;
assign R10C37_E26 = R10C37_Q6;
assign R10C37_W25 = R10C37_Q5;
assign R10C37_W26 = R10C37_Q6;
assign R10C37_E24 = R10C37_Q4;
assign R10C37_E27 = R10C37_Q7;
assign R10C37_W24 = R10C37_Q4;
assign R10C37_W27 = R10C37_Q7;
assign R10C37_E20 = R10C37_Q0;
assign R10C37_E23 = R10C37_Q3;
assign R10C37_W20 = R10C37_Q0;
assign R10C37_W23 = R10C37_Q3;
assign R10C37_B0 = R10C37_F3;
assign R10C37_B1 = R10C37_F3;
assign R10C37_B2 = R10C37_F1;
assign R10C37_B3 = R10C37_F1;
assign R10C37_B4 = R10C37_F1;
assign R10C37_B5 = R10C37_F1;
assign R10C37_B6 = R10C37_F1;
assign R10C37_B7 = R10C37_F1;
assign R10C37_D0 = R10C37_F2;
assign R10C37_D1 = R10C37_F2;
assign R10C37_D2 = R10C37_F0;
assign R10C37_D3 = R10C37_F0;
assign R10C37_D4 = R10C37_F0;
assign R10C37_D5 = R10C37_F0;
assign R10C37_D6 = R10C37_F0;
assign R10C37_D7 = R10C37_F0;
assign R10C37_X02 = R10C37_Q1;
assign R10C37_X04 = R10C37_Q7;
assign R10C37_X06 = R10C37_Q1;
assign R10C37_X08 = R10C37_Q7;
assign R10C37_X01 = R10C37_Q0;
assign R10C37_X03 = R10C37_Q6;
assign R10C37_X05 = R10C37_Q0;
assign R10C37_X07 = R10C37_Q6;
assign R10C37_N10 = R10C37_Q0;
assign R10C37_SN10 = R10C37_Q0;
assign R10C37_SN20 = R10C37_Q0;
assign R10C37_N13 = R10C37_Q0;
assign R10C37_S10 = R10C37_Q0;
assign R10C37_S13 = R10C37_Q0;
assign R10C37_E10 = R10C37_Q0;
assign R10C37_EW10 = R10C37_Q0;
assign R10C37_EW20 = R10C37_Q0;
assign R10C37_E13 = R10C37_Q0;
assign R10C37_W10 = R10C37_Q0;
assign R10C37_W13 = R10C37_Q0;
assign R10C37_E11 = R10C37_EW10;
assign R10C37_W11 = R10C37_EW10;
assign R10C37_E12 = R10C37_EW20;
assign R10C37_W12 = R10C37_EW20;
assign R10C37_S11 = R10C37_SN10;
assign R10C37_N11 = R10C37_SN10;
assign R10C37_S12 = R10C37_SN20;
assign R10C37_N12 = R10C37_SN20;
assign R10C40_CLK0 = VCC;
assign R10C40_CLK1 = VCC;
assign R10C40_CLK2 = VCC;
assign R10C40_LSR0 = VCC;
assign R10C40_LSR1 = VCC;
assign R10C40_LSR2 = VCC;
assign R10C40_CE0 = VCC;
assign R10C40_CE1 = VCC;
assign R10C40_CE2 = VCC;
assign R10C40_SEL0 = VCC;
assign R10C40_SEL1 = VCC;
assign R10C40_SEL2 = VCC;
assign R10C40_SEL3 = VCC;
assign R10C40_SEL4 = VCC;
assign R10C40_SEL5 = VCC;
assign R10C40_SEL6 = VCC;
assign R10C40_SEL7 = VCC;
assign R10C40_C0 = R10C40_F4;
assign R10C40_C1 = R10C40_F4;
assign R10C40_C2 = R10C40_F4;
assign R10C40_C3 = R10C40_F4;
assign R10C40_A4 = R10C40_F7;
assign R10C40_A5 = R10C40_F7;
assign R10C40_A6 = R10C40_F5;
assign R10C40_A7 = R10C40_F5;
assign R10C40_N82 = R10C40_Q4;
assign R10C40_S82 = R10C40_Q4;
assign R10C40_E82 = R10C40_Q4;
assign R10C40_W82 = R10C40_Q4;
assign R10C40_A0 = R10C40_F5;
assign R10C40_A1 = R10C40_F5;
assign R10C40_A2 = R10C40_F5;
assign R10C40_A3 = R10C40_F5;
assign R10C40_C4 = R10C40_F6;
assign R10C40_C5 = R10C40_F6;
assign R10C40_C6 = R10C40_F4;
assign R10C40_C7 = R10C40_F4;
assign R10C40_N81 = R10C40_Q1;
assign R10C40_S81 = R10C40_Q1;
assign R10C40_E81 = R10C40_Q1;
assign R10C40_W81 = R10C40_Q1;
assign R10C40_N21 = R10C40_Q1;
assign R10C40_N22 = R10C40_Q2;
assign R10C40_S21 = R10C40_Q1;
assign R10C40_S22 = R10C40_Q2;
assign R10C40_E21 = R10C40_Q1;
assign R10C40_E22 = R10C40_Q2;
assign R10C40_W21 = R10C40_Q1;
assign R10C40_W22 = R10C40_Q2;
assign R10C40_E80 = R10C40_Q0;
assign R10C40_W80 = R10C40_Q0;
assign R10C40_N25 = R10C40_Q5;
assign R10C40_N26 = R10C40_Q6;
assign R10C40_S25 = R10C40_Q5;
assign R10C40_S26 = R10C40_Q6;
assign R10C40_N83 = R10C40_Q5;
assign R10C40_S83 = R10C40_Q5;
assign R10C40_N24 = R10C40_Q4;
assign R10C40_N27 = R10C40_Q7;
assign R10C40_S24 = R10C40_Q4;
assign R10C40_S27 = R10C40_Q7;
assign R10C40_N20 = R10C40_Q0;
assign R10C40_N23 = R10C40_Q3;
assign R10C40_S20 = R10C40_Q0;
assign R10C40_S23 = R10C40_Q3;
assign R10C40_N80 = R10C40_Q0;
assign R10C40_S80 = R10C40_Q0;
assign R10C40_E83 = R10C40_Q5;
assign R10C40_W83 = R10C40_Q5;
assign R10C40_E25 = R10C40_Q5;
assign R10C40_E26 = R10C40_Q6;
assign R10C40_W25 = R10C40_Q5;
assign R10C40_W26 = R10C40_Q6;
assign R10C40_E24 = R10C40_Q4;
assign R10C40_E27 = R10C40_Q7;
assign R10C40_W24 = R10C40_Q4;
assign R10C40_W27 = R10C40_Q7;
assign R10C40_E20 = R10C40_Q0;
assign R10C40_E23 = R10C40_Q3;
assign R10C40_W20 = R10C40_Q0;
assign R10C40_W23 = R10C40_Q3;
assign R10C40_B0 = R10C40_F3;
assign R10C40_B1 = R10C40_F3;
assign R10C40_B2 = R10C40_F1;
assign R10C40_B3 = R10C40_F1;
assign R10C40_B4 = R10C40_F1;
assign R10C40_B5 = R10C40_F1;
assign R10C40_B6 = R10C40_F1;
assign R10C40_B7 = R10C40_F1;
assign R10C40_D0 = R10C40_F2;
assign R10C40_D1 = R10C40_F2;
assign R10C40_D2 = R10C40_F0;
assign R10C40_D3 = R10C40_F0;
assign R10C40_D4 = R10C40_F0;
assign R10C40_D5 = R10C40_F0;
assign R10C40_D6 = R10C40_F0;
assign R10C40_D7 = R10C40_F0;
assign R10C40_X02 = R10C40_Q1;
assign R10C40_X04 = R10C40_Q7;
assign R10C40_X06 = R10C40_Q1;
assign R10C40_X08 = R10C40_Q7;
assign R10C40_X01 = R10C40_Q0;
assign R10C40_X03 = R10C40_Q6;
assign R10C40_X05 = R10C40_Q0;
assign R10C40_X07 = R10C40_Q6;
assign R10C40_N10 = R10C40_Q0;
assign R10C40_SN10 = R10C40_Q0;
assign R10C40_SN20 = R10C40_Q0;
assign R10C40_N13 = R10C40_Q0;
assign R10C40_S10 = R10C40_Q0;
assign R10C40_S13 = R10C40_Q0;
assign R10C40_E10 = R10C40_Q0;
assign R10C40_EW10 = R10C40_Q0;
assign R10C40_EW20 = R10C40_Q0;
assign R10C40_E13 = R10C40_Q0;
assign R10C40_W10 = R10C40_Q0;
assign R10C40_W13 = R10C40_Q0;
assign R10C40_E11 = R10C40_EW10;
assign R10C40_W11 = R10C40_EW10;
assign R10C40_E12 = R10C40_EW20;
assign R10C40_W12 = R10C40_EW20;
assign R10C40_S11 = R10C40_SN10;
assign R10C40_N11 = R10C40_SN10;
assign R10C40_S12 = R10C40_SN20;
assign R10C40_N12 = R10C40_SN20;
assign R10C43_CLK0 = VCC;
assign R10C43_CLK1 = VCC;
assign R10C43_CLK2 = VCC;
assign R10C43_LSR0 = VCC;
assign R10C43_LSR1 = VCC;
assign R10C43_LSR2 = VCC;
assign R10C43_CE0 = VCC;
assign R10C43_CE1 = VCC;
assign R10C43_CE2 = VCC;
assign R10C43_SEL0 = VCC;
assign R10C43_SEL1 = VCC;
assign R10C43_SEL2 = VCC;
assign R10C43_SEL3 = VCC;
assign R10C43_SEL4 = VCC;
assign R10C43_SEL5 = VCC;
assign R10C43_SEL6 = VCC;
assign R10C43_SEL7 = VCC;
assign R10C43_C0 = R10C43_F4;
assign R10C43_C1 = R10C43_F4;
assign R10C43_C2 = R10C43_F4;
assign R10C43_C3 = R10C43_F4;
assign R10C43_A4 = R10C43_F7;
assign R10C43_A5 = R10C43_F7;
assign R10C43_A6 = R10C43_F5;
assign R10C43_A7 = R10C43_F5;
assign R10C43_N82 = R10C43_Q4;
assign R10C43_S82 = R10C43_Q4;
assign R10C43_E82 = R10C43_Q4;
assign R10C43_W82 = R10C43_Q4;
assign R10C43_A0 = R10C43_F5;
assign R10C43_A1 = R10C43_F5;
assign R10C43_A2 = R10C43_F5;
assign R10C43_A3 = R10C43_F5;
assign R10C43_C4 = R10C43_F6;
assign R10C43_C5 = R10C43_F6;
assign R10C43_C6 = R10C43_F4;
assign R10C43_C7 = R10C43_F4;
assign R10C43_N81 = R10C43_Q1;
assign R10C43_S81 = R10C43_Q1;
assign R10C43_E81 = R10C43_Q1;
assign R10C43_W81 = R10C43_Q1;
assign R10C43_N21 = R10C43_Q1;
assign R10C43_N22 = R10C43_Q2;
assign R10C43_S21 = R10C43_Q1;
assign R10C43_S22 = R10C43_Q2;
assign R10C43_E21 = R10C43_Q1;
assign R10C43_E22 = R10C43_Q2;
assign R10C43_W21 = R10C43_Q1;
assign R10C43_W22 = R10C43_Q2;
assign R10C43_E80 = R10C43_Q0;
assign R10C43_W80 = R10C43_Q0;
assign R10C43_N25 = R10C43_Q5;
assign R10C43_N26 = R10C43_Q6;
assign R10C43_S25 = R10C43_Q5;
assign R10C43_S26 = R10C43_Q6;
assign R10C43_N83 = R10C43_Q5;
assign R10C43_S83 = R10C43_Q5;
assign R10C43_N24 = R10C43_Q4;
assign R10C43_N27 = R10C43_Q7;
assign R10C43_S24 = R10C43_Q4;
assign R10C43_S27 = R10C43_Q7;
assign R10C43_N20 = R10C43_Q0;
assign R10C43_N23 = R10C43_Q3;
assign R10C43_S20 = R10C43_Q0;
assign R10C43_S23 = R10C43_Q3;
assign R10C43_N80 = R10C43_Q0;
assign R10C43_S80 = R10C43_Q0;
assign R10C43_E83 = R10C43_Q5;
assign R10C43_W83 = R10C43_Q5;
assign R10C43_E25 = R10C43_Q5;
assign R10C43_E26 = R10C43_Q6;
assign R10C43_W25 = R10C43_Q5;
assign R10C43_W26 = R10C43_Q6;
assign R10C43_E24 = R10C43_Q4;
assign R10C43_E27 = R10C43_Q7;
assign R10C43_W24 = R10C43_Q4;
assign R10C43_W27 = R10C43_Q7;
assign R10C43_E20 = R10C43_Q0;
assign R10C43_E23 = R10C43_Q3;
assign R10C43_W20 = R10C43_Q0;
assign R10C43_W23 = R10C43_Q3;
assign R10C43_B0 = R10C43_F3;
assign R10C43_B1 = R10C43_F3;
assign R10C43_B2 = R10C43_F1;
assign R10C43_B3 = R10C43_F1;
assign R10C43_B4 = R10C43_F1;
assign R10C43_B5 = R10C43_F1;
assign R10C43_B6 = R10C43_F1;
assign R10C43_B7 = R10C43_F1;
assign R10C43_D0 = R10C43_F2;
assign R10C43_D1 = R10C43_F2;
assign R10C43_D2 = R10C43_F0;
assign R10C43_D3 = R10C43_F0;
assign R10C43_D4 = R10C43_F0;
assign R10C43_D5 = R10C43_F0;
assign R10C43_D6 = R10C43_F0;
assign R10C43_D7 = R10C43_F0;
assign R10C43_X02 = R10C43_Q1;
assign R10C43_X04 = R10C43_Q7;
assign R10C43_X06 = R10C43_Q1;
assign R10C43_X08 = R10C43_Q7;
assign R10C43_X01 = R10C43_Q0;
assign R10C43_X03 = R10C43_Q6;
assign R10C43_X05 = R10C43_Q0;
assign R10C43_X07 = R10C43_Q6;
assign R10C43_N10 = R10C43_Q0;
assign R10C43_SN10 = R10C43_Q0;
assign R10C43_SN20 = R10C43_Q0;
assign R10C43_N13 = R10C43_Q0;
assign R10C43_S10 = R10C43_Q0;
assign R10C43_S13 = R10C43_Q0;
assign R10C43_E10 = R10C43_Q0;
assign R10C43_EW10 = R10C43_Q0;
assign R10C43_EW20 = R10C43_Q0;
assign R10C43_E13 = R10C43_Q0;
assign R10C43_W10 = R10C43_Q0;
assign R10C43_W13 = R10C43_Q0;
assign R10C43_E11 = R10C43_EW10;
assign R10C43_W11 = R10C43_EW10;
assign R10C43_E12 = R10C43_EW20;
assign R10C43_W12 = R10C43_EW20;
assign R10C43_S11 = R10C43_SN10;
assign R10C43_N11 = R10C43_SN10;
assign R10C43_S12 = R10C43_SN20;
assign R10C43_N12 = R10C43_SN20;
assign R28C4_CLK0 = VCC;
assign R28C4_CLK1 = VCC;
assign R28C4_CLK2 = VCC;
assign R28C4_LSR0 = VCC;
assign R28C4_LSR1 = VCC;
assign R28C4_LSR2 = VCC;
assign R28C4_CE0 = VCC;
assign R28C4_CE1 = VCC;
assign R28C4_CE2 = VCC;
assign R28C4_SEL0 = VCC;
assign R28C4_SEL1 = VCC;
assign R28C4_SEL2 = VCC;
assign R28C4_SEL3 = VCC;
assign R28C4_SEL4 = VCC;
assign R28C4_SEL5 = VCC;
assign R28C4_SEL6 = VCC;
assign R28C4_SEL7 = VCC;
assign R28C4_C0 = R28C4_F4;
assign R28C4_C1 = R28C4_F4;
assign R28C4_C2 = R28C4_F4;
assign R28C4_C3 = R28C4_F4;
assign R28C4_A4 = R28C4_F7;
assign R28C4_A5 = R28C4_F7;
assign R28C4_A6 = R28C4_F5;
assign R28C4_A7 = R28C4_F5;
assign R28C4_N82 = R28C4_Q4;
assign R28C4_S82 = R28C4_Q4;
assign R28C4_E82 = R28C4_Q4;
assign R28C4_W82 = R28C4_Q4;
assign R28C4_A0 = R28C4_F5;
assign R28C4_A1 = R28C4_F5;
assign R28C4_A2 = R28C4_F5;
assign R28C4_A3 = R28C4_F5;
assign R28C4_C4 = R28C4_F6;
assign R28C4_C5 = R28C4_F6;
assign R28C4_C6 = R28C4_F4;
assign R28C4_C7 = R28C4_F4;
assign R28C4_N81 = R28C4_Q1;
assign R28C4_S81 = R28C4_Q1;
assign R28C4_E81 = R28C4_Q1;
assign R28C4_W81 = R28C4_Q1;
assign R28C4_N21 = R28C4_Q1;
assign R28C4_N22 = R28C4_Q2;
assign R28C4_S21 = R28C4_Q1;
assign R28C4_S22 = R28C4_Q2;
assign R28C4_E21 = R28C4_Q1;
assign R28C4_E22 = R28C4_Q2;
assign R28C4_W21 = R28C4_Q1;
assign R28C4_W22 = R28C4_Q2;
assign R28C4_E80 = R28C4_Q0;
assign R28C4_W80 = R28C4_Q0;
assign R28C4_N25 = R28C4_Q5;
assign R28C4_N26 = R28C4_Q6;
assign R28C4_S25 = R28C4_Q5;
assign R28C4_S26 = R28C4_Q6;
assign R28C4_N83 = R28C4_Q5;
assign R28C4_S83 = R28C4_Q5;
assign R28C4_N24 = R28C4_Q4;
assign R28C4_N27 = R28C4_Q7;
assign R28C4_S24 = R28C4_Q4;
assign R28C4_S27 = R28C4_Q7;
assign R28C4_N20 = R28C4_Q0;
assign R28C4_N23 = R28C4_Q3;
assign R28C4_S20 = R28C4_Q0;
assign R28C4_S23 = R28C4_Q3;
assign R28C4_N80 = R28C4_Q0;
assign R28C4_S80 = R28C4_Q0;
assign R28C4_E83 = R28C4_Q5;
assign R28C4_W83 = R28C4_Q5;
assign R28C4_E25 = R28C4_Q5;
assign R28C4_E26 = R28C4_Q6;
assign R28C4_W25 = R28C4_Q5;
assign R28C4_W26 = R28C4_Q6;
assign R28C4_E24 = R28C4_Q4;
assign R28C4_E27 = R28C4_Q7;
assign R28C4_W24 = R28C4_Q4;
assign R28C4_W27 = R28C4_Q7;
assign R28C4_E20 = R28C4_Q0;
assign R28C4_E23 = R28C4_Q3;
assign R28C4_W20 = R28C4_Q0;
assign R28C4_W23 = R28C4_Q3;
assign R28C4_B0 = R28C4_F3;
assign R28C4_B1 = R28C4_F3;
assign R28C4_B2 = R28C4_F1;
assign R28C4_B3 = R28C4_F1;
assign R28C4_B4 = R28C4_F1;
assign R28C4_B5 = R28C4_F1;
assign R28C4_B6 = R28C4_F1;
assign R28C4_B7 = R28C4_F1;
assign R28C4_D0 = R28C4_F2;
assign R28C4_D1 = R28C4_F2;
assign R28C4_D2 = R28C4_F0;
assign R28C4_D3 = R28C4_F0;
assign R28C4_D4 = R28C4_F0;
assign R28C4_D5 = R28C4_F0;
assign R28C4_D6 = R28C4_F0;
assign R28C4_D7 = R28C4_F0;
assign R28C4_X02 = R28C4_Q1;
assign R28C4_X04 = R28C4_Q7;
assign R28C4_X06 = R28C4_Q1;
assign R28C4_X08 = R28C4_Q7;
assign R28C4_X01 = R28C4_Q0;
assign R28C4_X03 = R28C4_Q6;
assign R28C4_X05 = R28C4_Q0;
assign R28C4_X07 = R28C4_Q6;
assign R28C4_N10 = R28C4_Q0;
assign R28C4_SN10 = R28C4_Q0;
assign R28C4_SN20 = R28C4_Q0;
assign R28C4_N13 = R28C4_Q0;
assign R28C4_S10 = R28C4_Q0;
assign R28C4_S13 = R28C4_Q0;
assign R28C4_E10 = R28C4_Q0;
assign R28C4_EW10 = R28C4_Q0;
assign R28C4_EW20 = R28C4_Q0;
assign R28C4_E13 = R28C4_Q0;
assign R28C4_W10 = R28C4_Q0;
assign R28C4_W13 = R28C4_Q0;
assign R28C4_E11 = R28C4_EW10;
assign R28C4_W11 = R28C4_EW10;
assign R28C4_E12 = R28C4_EW20;
assign R28C4_W12 = R28C4_EW20;
assign R28C4_S11 = R28C4_SN10;
assign R28C4_N11 = R28C4_SN10;
assign R28C4_S12 = R28C4_SN20;
assign R28C4_N12 = R28C4_SN20;
assign R28C7_CLK0 = VCC;
assign R28C7_CLK1 = VCC;
assign R28C7_CLK2 = VCC;
assign R28C7_LSR0 = VCC;
assign R28C7_LSR1 = VCC;
assign R28C7_LSR2 = VCC;
assign R28C7_CE0 = VCC;
assign R28C7_CE1 = VCC;
assign R28C7_CE2 = VCC;
assign R28C7_SEL0 = VCC;
assign R28C7_SEL1 = VCC;
assign R28C7_SEL2 = VCC;
assign R28C7_SEL3 = VCC;
assign R28C7_SEL4 = VCC;
assign R28C7_SEL5 = VCC;
assign R28C7_SEL6 = VCC;
assign R28C7_SEL7 = VCC;
assign R28C7_C0 = R28C7_F4;
assign R28C7_C1 = R28C7_F4;
assign R28C7_C2 = R28C7_F4;
assign R28C7_C3 = R28C7_F4;
assign R28C7_A4 = R28C7_F7;
assign R28C7_A5 = R28C7_F7;
assign R28C7_A6 = R28C7_F5;
assign R28C7_A7 = R28C7_F5;
assign R28C7_N82 = R28C7_Q4;
assign R28C7_S82 = R28C7_Q4;
assign R28C7_E82 = R28C7_Q4;
assign R28C7_W82 = R28C7_Q4;
assign R28C7_A0 = R28C7_F5;
assign R28C7_A1 = R28C7_F5;
assign R28C7_A2 = R28C7_F5;
assign R28C7_A3 = R28C7_F5;
assign R28C7_C4 = R28C7_F6;
assign R28C7_C5 = R28C7_F6;
assign R28C7_C6 = R28C7_F4;
assign R28C7_C7 = R28C7_F4;
assign R28C7_N81 = R28C7_Q1;
assign R28C7_S81 = R28C7_Q1;
assign R28C7_E81 = R28C7_Q1;
assign R28C7_W81 = R28C7_Q1;
assign R28C7_N21 = R28C7_Q1;
assign R28C7_N22 = R28C7_Q2;
assign R28C7_S21 = R28C7_Q1;
assign R28C7_S22 = R28C7_Q2;
assign R28C7_E21 = R28C7_Q1;
assign R28C7_E22 = R28C7_Q2;
assign R28C7_W21 = R28C7_Q1;
assign R28C7_W22 = R28C7_Q2;
assign R28C7_E80 = R28C7_Q0;
assign R28C7_W80 = R28C7_Q0;
assign R28C7_N25 = R28C7_Q5;
assign R28C7_N26 = R28C7_Q6;
assign R28C7_S25 = R28C7_Q5;
assign R28C7_S26 = R28C7_Q6;
assign R28C7_N83 = R28C7_Q5;
assign R28C7_S83 = R28C7_Q5;
assign R28C7_N24 = R28C7_Q4;
assign R28C7_N27 = R28C7_Q7;
assign R28C7_S24 = R28C7_Q4;
assign R28C7_S27 = R28C7_Q7;
assign R28C7_N20 = R28C7_Q0;
assign R28C7_N23 = R28C7_Q3;
assign R28C7_S20 = R28C7_Q0;
assign R28C7_S23 = R28C7_Q3;
assign R28C7_N80 = R28C7_Q0;
assign R28C7_S80 = R28C7_Q0;
assign R28C7_E83 = R28C7_Q5;
assign R28C7_W83 = R28C7_Q5;
assign R28C7_E25 = R28C7_Q5;
assign R28C7_E26 = R28C7_Q6;
assign R28C7_W25 = R28C7_Q5;
assign R28C7_W26 = R28C7_Q6;
assign R28C7_E24 = R28C7_Q4;
assign R28C7_E27 = R28C7_Q7;
assign R28C7_W24 = R28C7_Q4;
assign R28C7_W27 = R28C7_Q7;
assign R28C7_E20 = R28C7_Q0;
assign R28C7_E23 = R28C7_Q3;
assign R28C7_W20 = R28C7_Q0;
assign R28C7_W23 = R28C7_Q3;
assign R28C7_B0 = R28C7_F3;
assign R28C7_B1 = R28C7_F3;
assign R28C7_B2 = R28C7_F1;
assign R28C7_B3 = R28C7_F1;
assign R28C7_B4 = R28C7_F1;
assign R28C7_B5 = R28C7_F1;
assign R28C7_B6 = R28C7_F1;
assign R28C7_B7 = R28C7_F1;
assign R28C7_D0 = R28C7_F2;
assign R28C7_D1 = R28C7_F2;
assign R28C7_D2 = R28C7_F0;
assign R28C7_D3 = R28C7_F0;
assign R28C7_D4 = R28C7_F0;
assign R28C7_D5 = R28C7_F0;
assign R28C7_D6 = R28C7_F0;
assign R28C7_D7 = R28C7_F0;
assign R28C7_X02 = R28C7_Q1;
assign R28C7_X04 = R28C7_Q7;
assign R28C7_X06 = R28C7_Q1;
assign R28C7_X08 = R28C7_Q7;
assign R28C7_X01 = R28C7_Q0;
assign R28C7_X03 = R28C7_Q6;
assign R28C7_X05 = R28C7_Q0;
assign R28C7_X07 = R28C7_Q6;
assign R28C7_N10 = R28C7_Q0;
assign R28C7_SN10 = R28C7_Q0;
assign R28C7_SN20 = R28C7_Q0;
assign R28C7_N13 = R28C7_Q0;
assign R28C7_S10 = R28C7_Q0;
assign R28C7_S13 = R28C7_Q0;
assign R28C7_E10 = R28C7_Q0;
assign R28C7_EW10 = R28C7_Q0;
assign R28C7_EW20 = R28C7_Q0;
assign R28C7_E13 = R28C7_Q0;
assign R28C7_W10 = R28C7_Q0;
assign R28C7_W13 = R28C7_Q0;
assign R28C7_E11 = R28C7_EW10;
assign R28C7_W11 = R28C7_EW10;
assign R28C7_E12 = R28C7_EW20;
assign R28C7_W12 = R28C7_EW20;
assign R28C7_S11 = R28C7_SN10;
assign R28C7_N11 = R28C7_SN10;
assign R28C7_S12 = R28C7_SN20;
assign R28C7_N12 = R28C7_SN20;
assign R28C10_CLK0 = VCC;
assign R28C10_CLK1 = VCC;
assign R28C10_CLK2 = VCC;
assign R28C10_LSR0 = VCC;
assign R28C10_LSR1 = VCC;
assign R28C10_LSR2 = VCC;
assign R28C10_CE0 = VCC;
assign R28C10_CE1 = VCC;
assign R28C10_CE2 = VCC;
assign R28C10_SEL0 = VCC;
assign R28C10_SEL1 = VCC;
assign R28C10_SEL2 = VCC;
assign R28C10_SEL3 = VCC;
assign R28C10_SEL4 = VCC;
assign R28C10_SEL5 = VCC;
assign R28C10_SEL6 = VCC;
assign R28C10_SEL7 = VCC;
assign R28C10_C0 = R28C10_F4;
assign R28C10_C1 = R28C10_F4;
assign R28C10_C2 = R28C10_F4;
assign R28C10_C3 = R28C10_F4;
assign R28C10_A4 = R28C10_F7;
assign R28C10_A5 = R28C10_F7;
assign R28C10_A6 = R28C10_F5;
assign R28C10_A7 = R28C10_F5;
assign R28C10_N82 = R28C10_Q4;
assign R28C10_S82 = R28C10_Q4;
assign R28C10_E82 = R28C10_Q4;
assign R28C10_W82 = R28C10_Q4;
assign R28C10_A0 = R28C10_F5;
assign R28C10_A1 = R28C10_F5;
assign R28C10_A2 = R28C10_F5;
assign R28C10_A3 = R28C10_F5;
assign R28C10_C4 = R28C10_F6;
assign R28C10_C5 = R28C10_F6;
assign R28C10_C6 = R28C10_F4;
assign R28C10_C7 = R28C10_F4;
assign R28C10_N81 = R28C10_Q1;
assign R28C10_S81 = R28C10_Q1;
assign R28C10_E81 = R28C10_Q1;
assign R28C10_W81 = R28C10_Q1;
assign R28C10_N21 = R28C10_Q1;
assign R28C10_N22 = R28C10_Q2;
assign R28C10_S21 = R28C10_Q1;
assign R28C10_S22 = R28C10_Q2;
assign R28C10_E21 = R28C10_Q1;
assign R28C10_E22 = R28C10_Q2;
assign R28C10_W21 = R28C10_Q1;
assign R28C10_W22 = R28C10_Q2;
assign R28C10_E80 = R28C10_Q0;
assign R28C10_W80 = R28C10_Q0;
assign R28C10_N25 = R28C10_Q5;
assign R28C10_N26 = R28C10_Q6;
assign R28C10_S25 = R28C10_Q5;
assign R28C10_S26 = R28C10_Q6;
assign R28C10_N83 = R28C10_Q5;
assign R28C10_S83 = R28C10_Q5;
assign R28C10_N24 = R28C10_Q4;
assign R28C10_N27 = R28C10_Q7;
assign R28C10_S24 = R28C10_Q4;
assign R28C10_S27 = R28C10_Q7;
assign R28C10_N20 = R28C10_Q0;
assign R28C10_N23 = R28C10_Q3;
assign R28C10_S20 = R28C10_Q0;
assign R28C10_S23 = R28C10_Q3;
assign R28C10_N80 = R28C10_Q0;
assign R28C10_S80 = R28C10_Q0;
assign R28C10_E83 = R28C10_Q5;
assign R28C10_W83 = R28C10_Q5;
assign R28C10_E25 = R28C10_Q5;
assign R28C10_E26 = R28C10_Q6;
assign R28C10_W25 = R28C10_Q5;
assign R28C10_W26 = R28C10_Q6;
assign R28C10_E24 = R28C10_Q4;
assign R28C10_E27 = R28C10_Q7;
assign R28C10_W24 = R28C10_Q4;
assign R28C10_W27 = R28C10_Q7;
assign R28C10_E20 = R28C10_Q0;
assign R28C10_E23 = R28C10_Q3;
assign R28C10_W20 = R28C10_Q0;
assign R28C10_W23 = R28C10_Q3;
assign R28C10_B0 = R28C10_F3;
assign R28C10_B1 = R28C10_F3;
assign R28C10_B2 = R28C10_F1;
assign R28C10_B3 = R28C10_F1;
assign R28C10_B4 = R28C10_F1;
assign R28C10_B5 = R28C10_F1;
assign R28C10_B6 = R28C10_F1;
assign R28C10_B7 = R28C10_F1;
assign R28C10_D0 = R28C10_F2;
assign R28C10_D1 = R28C10_F2;
assign R28C10_D2 = R28C10_F0;
assign R28C10_D3 = R28C10_F0;
assign R28C10_D4 = R28C10_F0;
assign R28C10_D5 = R28C10_F0;
assign R28C10_D6 = R28C10_F0;
assign R28C10_D7 = R28C10_F0;
assign R28C10_X02 = R28C10_Q1;
assign R28C10_X04 = R28C10_Q7;
assign R28C10_X06 = R28C10_Q1;
assign R28C10_X08 = R28C10_Q7;
assign R28C10_X01 = R28C10_Q0;
assign R28C10_X03 = R28C10_Q6;
assign R28C10_X05 = R28C10_Q0;
assign R28C10_X07 = R28C10_Q6;
assign R28C10_N10 = R28C10_Q0;
assign R28C10_SN10 = R28C10_Q0;
assign R28C10_SN20 = R28C10_Q0;
assign R28C10_N13 = R28C10_Q0;
assign R28C10_S10 = R28C10_Q0;
assign R28C10_S13 = R28C10_Q0;
assign R28C10_E10 = R28C10_Q0;
assign R28C10_EW10 = R28C10_Q0;
assign R28C10_EW20 = R28C10_Q0;
assign R28C10_E13 = R28C10_Q0;
assign R28C10_W10 = R28C10_Q0;
assign R28C10_W13 = R28C10_Q0;
assign R28C10_E11 = R28C10_EW10;
assign R28C10_W11 = R28C10_EW10;
assign R28C10_E12 = R28C10_EW20;
assign R28C10_W12 = R28C10_EW20;
assign R28C10_S11 = R28C10_SN10;
assign R28C10_N11 = R28C10_SN10;
assign R28C10_S12 = R28C10_SN20;
assign R28C10_N12 = R28C10_SN20;
assign R28C13_CLK0 = VCC;
assign R28C13_CLK1 = VCC;
assign R28C13_CLK2 = VCC;
assign R28C13_LSR0 = VCC;
assign R28C13_LSR1 = VCC;
assign R28C13_LSR2 = VCC;
assign R28C13_CE0 = VCC;
assign R28C13_CE1 = VCC;
assign R28C13_CE2 = VCC;
assign R28C13_SEL0 = VCC;
assign R28C13_SEL1 = VCC;
assign R28C13_SEL2 = VCC;
assign R28C13_SEL3 = VCC;
assign R28C13_SEL4 = VCC;
assign R28C13_SEL5 = VCC;
assign R28C13_SEL6 = VCC;
assign R28C13_SEL7 = VCC;
assign R28C13_C0 = R28C13_F4;
assign R28C13_C1 = R28C13_F4;
assign R28C13_C2 = R28C13_F4;
assign R28C13_C3 = R28C13_F4;
assign R28C13_A4 = R28C13_F7;
assign R28C13_A5 = R28C13_F7;
assign R28C13_A6 = R28C13_F5;
assign R28C13_A7 = R28C13_F5;
assign R28C13_N82 = R28C13_Q4;
assign R28C13_S82 = R28C13_Q4;
assign R28C13_E82 = R28C13_Q4;
assign R28C13_W82 = R28C13_Q4;
assign R28C13_A0 = R28C13_F5;
assign R28C13_A1 = R28C13_F5;
assign R28C13_A2 = R28C13_F5;
assign R28C13_A3 = R28C13_F5;
assign R28C13_C4 = R28C13_F6;
assign R28C13_C5 = R28C13_F6;
assign R28C13_C6 = R28C13_F4;
assign R28C13_C7 = R28C13_F4;
assign R28C13_N81 = R28C13_Q1;
assign R28C13_S81 = R28C13_Q1;
assign R28C13_E81 = R28C13_Q1;
assign R28C13_W81 = R28C13_Q1;
assign R28C13_N21 = R28C13_Q1;
assign R28C13_N22 = R28C13_Q2;
assign R28C13_S21 = R28C13_Q1;
assign R28C13_S22 = R28C13_Q2;
assign R28C13_E21 = R28C13_Q1;
assign R28C13_E22 = R28C13_Q2;
assign R28C13_W21 = R28C13_Q1;
assign R28C13_W22 = R28C13_Q2;
assign R28C13_E80 = R28C13_Q0;
assign R28C13_W80 = R28C13_Q0;
assign R28C13_N25 = R28C13_Q5;
assign R28C13_N26 = R28C13_Q6;
assign R28C13_S25 = R28C13_Q5;
assign R28C13_S26 = R28C13_Q6;
assign R28C13_N83 = R28C13_Q5;
assign R28C13_S83 = R28C13_Q5;
assign R28C13_N24 = R28C13_Q4;
assign R28C13_N27 = R28C13_Q7;
assign R28C13_S24 = R28C13_Q4;
assign R28C13_S27 = R28C13_Q7;
assign R28C13_N20 = R28C13_Q0;
assign R28C13_N23 = R28C13_Q3;
assign R28C13_S20 = R28C13_Q0;
assign R28C13_S23 = R28C13_Q3;
assign R28C13_N80 = R28C13_Q0;
assign R28C13_S80 = R28C13_Q0;
assign R28C13_E83 = R28C13_Q5;
assign R28C13_W83 = R28C13_Q5;
assign R28C13_E25 = R28C13_Q5;
assign R28C13_E26 = R28C13_Q6;
assign R28C13_W25 = R28C13_Q5;
assign R28C13_W26 = R28C13_Q6;
assign R28C13_E24 = R28C13_Q4;
assign R28C13_E27 = R28C13_Q7;
assign R28C13_W24 = R28C13_Q4;
assign R28C13_W27 = R28C13_Q7;
assign R28C13_E20 = R28C13_Q0;
assign R28C13_E23 = R28C13_Q3;
assign R28C13_W20 = R28C13_Q0;
assign R28C13_W23 = R28C13_Q3;
assign R28C13_B0 = R28C13_F3;
assign R28C13_B1 = R28C13_F3;
assign R28C13_B2 = R28C13_F1;
assign R28C13_B3 = R28C13_F1;
assign R28C13_B4 = R28C13_F1;
assign R28C13_B5 = R28C13_F1;
assign R28C13_B6 = R28C13_F1;
assign R28C13_B7 = R28C13_F1;
assign R28C13_D0 = R28C13_F2;
assign R28C13_D1 = R28C13_F2;
assign R28C13_D2 = R28C13_F0;
assign R28C13_D3 = R28C13_F0;
assign R28C13_D4 = R28C13_F0;
assign R28C13_D5 = R28C13_F0;
assign R28C13_D6 = R28C13_F0;
assign R28C13_D7 = R28C13_F0;
assign R28C13_X02 = R28C13_Q1;
assign R28C13_X04 = R28C13_Q7;
assign R28C13_X06 = R28C13_Q1;
assign R28C13_X08 = R28C13_Q7;
assign R28C13_X01 = R28C13_Q0;
assign R28C13_X03 = R28C13_Q6;
assign R28C13_X05 = R28C13_Q0;
assign R28C13_X07 = R28C13_Q6;
assign R28C13_N10 = R28C13_Q0;
assign R28C13_SN10 = R28C13_Q0;
assign R28C13_SN20 = R28C13_Q0;
assign R28C13_N13 = R28C13_Q0;
assign R28C13_S10 = R28C13_Q0;
assign R28C13_S13 = R28C13_Q0;
assign R28C13_E10 = R28C13_Q0;
assign R28C13_EW10 = R28C13_Q0;
assign R28C13_EW20 = R28C13_Q0;
assign R28C13_E13 = R28C13_Q0;
assign R28C13_W10 = R28C13_Q0;
assign R28C13_W13 = R28C13_Q0;
assign R28C13_E11 = R28C13_EW10;
assign R28C13_W11 = R28C13_EW10;
assign R28C13_E12 = R28C13_EW20;
assign R28C13_W12 = R28C13_EW20;
assign R28C13_S11 = R28C13_SN10;
assign R28C13_N11 = R28C13_SN10;
assign R28C13_S12 = R28C13_SN20;
assign R28C13_N12 = R28C13_SN20;
assign R28C16_CLK0 = VCC;
assign R28C16_CLK1 = VCC;
assign R28C16_CLK2 = VCC;
assign R28C16_LSR0 = VCC;
assign R28C16_LSR1 = VCC;
assign R28C16_LSR2 = VCC;
assign R28C16_CE0 = VCC;
assign R28C16_CE1 = VCC;
assign R28C16_CE2 = VCC;
assign R28C16_SEL0 = VCC;
assign R28C16_SEL1 = VCC;
assign R28C16_SEL2 = VCC;
assign R28C16_SEL3 = VCC;
assign R28C16_SEL4 = VCC;
assign R28C16_SEL5 = VCC;
assign R28C16_SEL6 = VCC;
assign R28C16_SEL7 = VCC;
assign R28C16_C0 = R28C16_F4;
assign R28C16_C1 = R28C16_F4;
assign R28C16_C2 = R28C16_F4;
assign R28C16_C3 = R28C16_F4;
assign R28C16_A4 = R28C16_F7;
assign R28C16_A5 = R28C16_F7;
assign R28C16_A6 = R28C16_F5;
assign R28C16_A7 = R28C16_F5;
assign R28C16_N82 = R28C16_Q4;
assign R28C16_S82 = R28C16_Q4;
assign R28C16_E82 = R28C16_Q4;
assign R28C16_W82 = R28C16_Q4;
assign R28C16_A0 = R28C16_F5;
assign R28C16_A1 = R28C16_F5;
assign R28C16_A2 = R28C16_F5;
assign R28C16_A3 = R28C16_F5;
assign R28C16_C4 = R28C16_F6;
assign R28C16_C5 = R28C16_F6;
assign R28C16_C6 = R28C16_F4;
assign R28C16_C7 = R28C16_F4;
assign R28C16_N81 = R28C16_Q1;
assign R28C16_S81 = R28C16_Q1;
assign R28C16_E81 = R28C16_Q1;
assign R28C16_W81 = R28C16_Q1;
assign R28C16_N21 = R28C16_Q1;
assign R28C16_N22 = R28C16_Q2;
assign R28C16_S21 = R28C16_Q1;
assign R28C16_S22 = R28C16_Q2;
assign R28C16_E21 = R28C16_Q1;
assign R28C16_E22 = R28C16_Q2;
assign R28C16_W21 = R28C16_Q1;
assign R28C16_W22 = R28C16_Q2;
assign R28C16_E80 = R28C16_Q0;
assign R28C16_W80 = R28C16_Q0;
assign R28C16_N25 = R28C16_Q5;
assign R28C16_N26 = R28C16_Q6;
assign R28C16_S25 = R28C16_Q5;
assign R28C16_S26 = R28C16_Q6;
assign R28C16_N83 = R28C16_Q5;
assign R28C16_S83 = R28C16_Q5;
assign R28C16_N24 = R28C16_Q4;
assign R28C16_N27 = R28C16_Q7;
assign R28C16_S24 = R28C16_Q4;
assign R28C16_S27 = R28C16_Q7;
assign R28C16_N20 = R28C16_Q0;
assign R28C16_N23 = R28C16_Q3;
assign R28C16_S20 = R28C16_Q0;
assign R28C16_S23 = R28C16_Q3;
assign R28C16_N80 = R28C16_Q0;
assign R28C16_S80 = R28C16_Q0;
assign R28C16_E83 = R28C16_Q5;
assign R28C16_W83 = R28C16_Q5;
assign R28C16_E25 = R28C16_Q5;
assign R28C16_E26 = R28C16_Q6;
assign R28C16_W25 = R28C16_Q5;
assign R28C16_W26 = R28C16_Q6;
assign R28C16_E24 = R28C16_Q4;
assign R28C16_E27 = R28C16_Q7;
assign R28C16_W24 = R28C16_Q4;
assign R28C16_W27 = R28C16_Q7;
assign R28C16_E20 = R28C16_Q0;
assign R28C16_E23 = R28C16_Q3;
assign R28C16_W20 = R28C16_Q0;
assign R28C16_W23 = R28C16_Q3;
assign R28C16_B0 = R28C16_F3;
assign R28C16_B1 = R28C16_F3;
assign R28C16_B2 = R28C16_F1;
assign R28C16_B3 = R28C16_F1;
assign R28C16_B4 = R28C16_F1;
assign R28C16_B5 = R28C16_F1;
assign R28C16_B6 = R28C16_F1;
assign R28C16_B7 = R28C16_F1;
assign R28C16_D0 = R28C16_F2;
assign R28C16_D1 = R28C16_F2;
assign R28C16_D2 = R28C16_F0;
assign R28C16_D3 = R28C16_F0;
assign R28C16_D4 = R28C16_F0;
assign R28C16_D5 = R28C16_F0;
assign R28C16_D6 = R28C16_F0;
assign R28C16_D7 = R28C16_F0;
assign R28C16_X02 = R28C16_Q1;
assign R28C16_X04 = R28C16_Q7;
assign R28C16_X06 = R28C16_Q1;
assign R28C16_X08 = R28C16_Q7;
assign R28C16_X01 = R28C16_Q0;
assign R28C16_X03 = R28C16_Q6;
assign R28C16_X05 = R28C16_Q0;
assign R28C16_X07 = R28C16_Q6;
assign R28C16_N10 = R28C16_Q0;
assign R28C16_SN10 = R28C16_Q0;
assign R28C16_SN20 = R28C16_Q0;
assign R28C16_N13 = R28C16_Q0;
assign R28C16_S10 = R28C16_Q0;
assign R28C16_S13 = R28C16_Q0;
assign R28C16_E10 = R28C16_Q0;
assign R28C16_EW10 = R28C16_Q0;
assign R28C16_EW20 = R28C16_Q0;
assign R28C16_E13 = R28C16_Q0;
assign R28C16_W10 = R28C16_Q0;
assign R28C16_W13 = R28C16_Q0;
assign R28C16_E11 = R28C16_EW10;
assign R28C16_W11 = R28C16_EW10;
assign R28C16_E12 = R28C16_EW20;
assign R28C16_W12 = R28C16_EW20;
assign R28C16_S11 = R28C16_SN10;
assign R28C16_N11 = R28C16_SN10;
assign R28C16_S12 = R28C16_SN20;
assign R28C16_N12 = R28C16_SN20;
assign R28C19_CLK0 = VCC;
assign R28C19_CLK1 = VCC;
assign R28C19_CLK2 = VCC;
assign R28C19_LSR0 = VCC;
assign R28C19_LSR1 = VCC;
assign R28C19_LSR2 = VCC;
assign R28C19_CE0 = VCC;
assign R28C19_CE1 = VCC;
assign R28C19_CE2 = VCC;
assign R28C19_SEL0 = VCC;
assign R28C19_SEL1 = VCC;
assign R28C19_SEL2 = VCC;
assign R28C19_SEL3 = VCC;
assign R28C19_SEL4 = VCC;
assign R28C19_SEL5 = VCC;
assign R28C19_SEL6 = VCC;
assign R28C19_SEL7 = VCC;
assign R28C19_C0 = R28C19_F4;
assign R28C19_C1 = R28C19_F4;
assign R28C19_C2 = R28C19_F4;
assign R28C19_C3 = R28C19_F4;
assign R28C19_A4 = R28C19_F7;
assign R28C19_A5 = R28C19_F7;
assign R28C19_A6 = R28C19_F5;
assign R28C19_A7 = R28C19_F5;
assign R28C19_N82 = R28C19_Q4;
assign R28C19_S82 = R28C19_Q4;
assign R28C19_E82 = R28C19_Q4;
assign R28C19_W82 = R28C19_Q4;
assign R28C19_A0 = R28C19_F5;
assign R28C19_A1 = R28C19_F5;
assign R28C19_A2 = R28C19_F5;
assign R28C19_A3 = R28C19_F5;
assign R28C19_C4 = R28C19_F6;
assign R28C19_C5 = R28C19_F6;
assign R28C19_C6 = R28C19_F4;
assign R28C19_C7 = R28C19_F4;
assign R28C19_N81 = R28C19_Q1;
assign R28C19_S81 = R28C19_Q1;
assign R28C19_E81 = R28C19_Q1;
assign R28C19_W81 = R28C19_Q1;
assign R28C19_N21 = R28C19_Q1;
assign R28C19_N22 = R28C19_Q2;
assign R28C19_S21 = R28C19_Q1;
assign R28C19_S22 = R28C19_Q2;
assign R28C19_E21 = R28C19_Q1;
assign R28C19_E22 = R28C19_Q2;
assign R28C19_W21 = R28C19_Q1;
assign R28C19_W22 = R28C19_Q2;
assign R28C19_E80 = R28C19_Q0;
assign R28C19_W80 = R28C19_Q0;
assign R28C19_N25 = R28C19_Q5;
assign R28C19_N26 = R28C19_Q6;
assign R28C19_S25 = R28C19_Q5;
assign R28C19_S26 = R28C19_Q6;
assign R28C19_N83 = R28C19_Q5;
assign R28C19_S83 = R28C19_Q5;
assign R28C19_N24 = R28C19_Q4;
assign R28C19_N27 = R28C19_Q7;
assign R28C19_S24 = R28C19_Q4;
assign R28C19_S27 = R28C19_Q7;
assign R28C19_N20 = R28C19_Q0;
assign R28C19_N23 = R28C19_Q3;
assign R28C19_S20 = R28C19_Q0;
assign R28C19_S23 = R28C19_Q3;
assign R28C19_N80 = R28C19_Q0;
assign R28C19_S80 = R28C19_Q0;
assign R28C19_E83 = R28C19_Q5;
assign R28C19_W83 = R28C19_Q5;
assign R28C19_E25 = R28C19_Q5;
assign R28C19_E26 = R28C19_Q6;
assign R28C19_W25 = R28C19_Q5;
assign R28C19_W26 = R28C19_Q6;
assign R28C19_E24 = R28C19_Q4;
assign R28C19_E27 = R28C19_Q7;
assign R28C19_W24 = R28C19_Q4;
assign R28C19_W27 = R28C19_Q7;
assign R28C19_E20 = R28C19_Q0;
assign R28C19_E23 = R28C19_Q3;
assign R28C19_W20 = R28C19_Q0;
assign R28C19_W23 = R28C19_Q3;
assign R28C19_B0 = R28C19_F3;
assign R28C19_B1 = R28C19_F3;
assign R28C19_B2 = R28C19_F1;
assign R28C19_B3 = R28C19_F1;
assign R28C19_B4 = R28C19_F1;
assign R28C19_B5 = R28C19_F1;
assign R28C19_B6 = R28C19_F1;
assign R28C19_B7 = R28C19_F1;
assign R28C19_D0 = R28C19_F2;
assign R28C19_D1 = R28C19_F2;
assign R28C19_D2 = R28C19_F0;
assign R28C19_D3 = R28C19_F0;
assign R28C19_D4 = R28C19_F0;
assign R28C19_D5 = R28C19_F0;
assign R28C19_D6 = R28C19_F0;
assign R28C19_D7 = R28C19_F0;
assign R28C19_X02 = R28C19_Q1;
assign R28C19_X04 = R28C19_Q7;
assign R28C19_X06 = R28C19_Q1;
assign R28C19_X08 = R28C19_Q7;
assign R28C19_X01 = R28C19_Q0;
assign R28C19_X03 = R28C19_Q6;
assign R28C19_X05 = R28C19_Q0;
assign R28C19_X07 = R28C19_Q6;
assign R28C19_N10 = R28C19_Q0;
assign R28C19_SN10 = R28C19_Q0;
assign R28C19_SN20 = R28C19_Q0;
assign R28C19_N13 = R28C19_Q0;
assign R28C19_S10 = R28C19_Q0;
assign R28C19_S13 = R28C19_Q0;
assign R28C19_E10 = R28C19_Q0;
assign R28C19_EW10 = R28C19_Q0;
assign R28C19_EW20 = R28C19_Q0;
assign R28C19_E13 = R28C19_Q0;
assign R28C19_W10 = R28C19_Q0;
assign R28C19_W13 = R28C19_Q0;
assign R28C19_E11 = R28C19_EW10;
assign R28C19_W11 = R28C19_EW10;
assign R28C19_E12 = R28C19_EW20;
assign R28C19_W12 = R28C19_EW20;
assign R28C19_S11 = R28C19_SN10;
assign R28C19_N11 = R28C19_SN10;
assign R28C19_S12 = R28C19_SN20;
assign R28C19_N12 = R28C19_SN20;
assign R28C22_CLK0 = VCC;
assign R28C22_CLK1 = VCC;
assign R28C22_CLK2 = VCC;
assign R28C22_LSR0 = VCC;
assign R28C22_LSR1 = VCC;
assign R28C22_LSR2 = VCC;
assign R28C22_CE0 = VCC;
assign R28C22_CE1 = VCC;
assign R28C22_CE2 = VCC;
assign R28C22_SEL0 = VCC;
assign R28C22_SEL1 = VCC;
assign R28C22_SEL2 = VCC;
assign R28C22_SEL3 = VCC;
assign R28C22_SEL4 = VCC;
assign R28C22_SEL5 = VCC;
assign R28C22_SEL6 = VCC;
assign R28C22_SEL7 = VCC;
assign R28C22_C0 = R28C22_F4;
assign R28C22_C1 = R28C22_F4;
assign R28C22_C2 = R28C22_F4;
assign R28C22_C3 = R28C22_F4;
assign R28C22_A4 = R28C22_F7;
assign R28C22_A5 = R28C22_F7;
assign R28C22_A6 = R28C22_F5;
assign R28C22_A7 = R28C22_F5;
assign R28C22_N82 = R28C22_Q4;
assign R28C22_S82 = R28C22_Q4;
assign R28C22_E82 = R28C22_Q4;
assign R28C22_W82 = R28C22_Q4;
assign R28C22_A0 = R28C22_F5;
assign R28C22_A1 = R28C22_F5;
assign R28C22_A2 = R28C22_F5;
assign R28C22_A3 = R28C22_F5;
assign R28C22_C4 = R28C22_F6;
assign R28C22_C5 = R28C22_F6;
assign R28C22_C6 = R28C22_F4;
assign R28C22_C7 = R28C22_F4;
assign R28C22_N81 = R28C22_Q1;
assign R28C22_S81 = R28C22_Q1;
assign R28C22_E81 = R28C22_Q1;
assign R28C22_W81 = R28C22_Q1;
assign R28C22_N21 = R28C22_Q1;
assign R28C22_N22 = R28C22_Q2;
assign R28C22_S21 = R28C22_Q1;
assign R28C22_S22 = R28C22_Q2;
assign R28C22_E21 = R28C22_Q1;
assign R28C22_E22 = R28C22_Q2;
assign R28C22_W21 = R28C22_Q1;
assign R28C22_W22 = R28C22_Q2;
assign R28C22_E80 = R28C22_Q0;
assign R28C22_W80 = R28C22_Q0;
assign R28C22_N25 = R28C22_Q5;
assign R28C22_N26 = R28C22_Q6;
assign R28C22_S25 = R28C22_Q5;
assign R28C22_S26 = R28C22_Q6;
assign R28C22_N83 = R28C22_Q5;
assign R28C22_S83 = R28C22_Q5;
assign R28C22_N24 = R28C22_Q4;
assign R28C22_N27 = R28C22_Q7;
assign R28C22_S24 = R28C22_Q4;
assign R28C22_S27 = R28C22_Q7;
assign R28C22_N20 = R28C22_Q0;
assign R28C22_N23 = R28C22_Q3;
assign R28C22_S20 = R28C22_Q0;
assign R28C22_S23 = R28C22_Q3;
assign R28C22_N80 = R28C22_Q0;
assign R28C22_S80 = R28C22_Q0;
assign R28C22_E83 = R28C22_Q5;
assign R28C22_W83 = R28C22_Q5;
assign R28C22_E25 = R28C22_Q5;
assign R28C22_E26 = R28C22_Q6;
assign R28C22_W25 = R28C22_Q5;
assign R28C22_W26 = R28C22_Q6;
assign R28C22_E24 = R28C22_Q4;
assign R28C22_E27 = R28C22_Q7;
assign R28C22_W24 = R28C22_Q4;
assign R28C22_W27 = R28C22_Q7;
assign R28C22_E20 = R28C22_Q0;
assign R28C22_E23 = R28C22_Q3;
assign R28C22_W20 = R28C22_Q0;
assign R28C22_W23 = R28C22_Q3;
assign R28C22_B0 = R28C22_F3;
assign R28C22_B1 = R28C22_F3;
assign R28C22_B2 = R28C22_F1;
assign R28C22_B3 = R28C22_F1;
assign R28C22_B4 = R28C22_F1;
assign R28C22_B5 = R28C22_F1;
assign R28C22_B6 = R28C22_F1;
assign R28C22_B7 = R28C22_F1;
assign R28C22_D0 = R28C22_F2;
assign R28C22_D1 = R28C22_F2;
assign R28C22_D2 = R28C22_F0;
assign R28C22_D3 = R28C22_F0;
assign R28C22_D4 = R28C22_F0;
assign R28C22_D5 = R28C22_F0;
assign R28C22_D6 = R28C22_F0;
assign R28C22_D7 = R28C22_F0;
assign R28C22_X02 = R28C22_Q1;
assign R28C22_X04 = R28C22_Q7;
assign R28C22_X06 = R28C22_Q1;
assign R28C22_X08 = R28C22_Q7;
assign R28C22_X01 = R28C22_Q0;
assign R28C22_X03 = R28C22_Q6;
assign R28C22_X05 = R28C22_Q0;
assign R28C22_X07 = R28C22_Q6;
assign R28C22_N10 = R28C22_Q0;
assign R28C22_SN10 = R28C22_Q0;
assign R28C22_SN20 = R28C22_Q0;
assign R28C22_N13 = R28C22_Q0;
assign R28C22_S10 = R28C22_Q0;
assign R28C22_S13 = R28C22_Q0;
assign R28C22_E10 = R28C22_Q0;
assign R28C22_EW10 = R28C22_Q0;
assign R28C22_EW20 = R28C22_Q0;
assign R28C22_E13 = R28C22_Q0;
assign R28C22_W10 = R28C22_Q0;
assign R28C22_W13 = R28C22_Q0;
assign R28C22_E11 = R28C22_EW10;
assign R28C22_W11 = R28C22_EW10;
assign R28C22_E12 = R28C22_EW20;
assign R28C22_W12 = R28C22_EW20;
assign R28C22_S11 = R28C22_SN10;
assign R28C22_N11 = R28C22_SN10;
assign R28C22_S12 = R28C22_SN20;
assign R28C22_N12 = R28C22_SN20;
assign R28C25_CLK0 = VCC;
assign R28C25_CLK1 = VCC;
assign R28C25_CLK2 = VCC;
assign R28C25_LSR0 = VCC;
assign R28C25_LSR1 = VCC;
assign R28C25_LSR2 = VCC;
assign R28C25_CE0 = VCC;
assign R28C25_CE1 = VCC;
assign R28C25_CE2 = VCC;
assign R28C25_SEL0 = VCC;
assign R28C25_SEL1 = VCC;
assign R28C25_SEL2 = VCC;
assign R28C25_SEL3 = VCC;
assign R28C25_SEL4 = VCC;
assign R28C25_SEL5 = VCC;
assign R28C25_SEL6 = VCC;
assign R28C25_SEL7 = VCC;
assign R28C25_C0 = R28C25_F4;
assign R28C25_C1 = R28C25_F4;
assign R28C25_C2 = R28C25_F4;
assign R28C25_C3 = R28C25_F4;
assign R28C25_A4 = R28C25_F7;
assign R28C25_A5 = R28C25_F7;
assign R28C25_A6 = R28C25_F5;
assign R28C25_A7 = R28C25_F5;
assign R28C25_N82 = R28C25_Q4;
assign R28C25_S82 = R28C25_Q4;
assign R28C25_E82 = R28C25_Q4;
assign R28C25_W82 = R28C25_Q4;
assign R28C25_A0 = R28C25_F5;
assign R28C25_A1 = R28C25_F5;
assign R28C25_A2 = R28C25_F5;
assign R28C25_A3 = R28C25_F5;
assign R28C25_C4 = R28C25_F6;
assign R28C25_C5 = R28C25_F6;
assign R28C25_C6 = R28C25_F4;
assign R28C25_C7 = R28C25_F4;
assign R28C25_N81 = R28C25_Q1;
assign R28C25_S81 = R28C25_Q1;
assign R28C25_E81 = R28C25_Q1;
assign R28C25_W81 = R28C25_Q1;
assign R28C25_N21 = R28C25_Q1;
assign R28C25_N22 = R28C25_Q2;
assign R28C25_S21 = R28C25_Q1;
assign R28C25_S22 = R28C25_Q2;
assign R28C25_E21 = R28C25_Q1;
assign R28C25_E22 = R28C25_Q2;
assign R28C25_W21 = R28C25_Q1;
assign R28C25_W22 = R28C25_Q2;
assign R28C25_E80 = R28C25_Q0;
assign R28C25_W80 = R28C25_Q0;
assign R28C25_N25 = R28C25_Q5;
assign R28C25_N26 = R28C25_Q6;
assign R28C25_S25 = R28C25_Q5;
assign R28C25_S26 = R28C25_Q6;
assign R28C25_N83 = R28C25_Q5;
assign R28C25_S83 = R28C25_Q5;
assign R28C25_N24 = R28C25_Q4;
assign R28C25_N27 = R28C25_Q7;
assign R28C25_S24 = R28C25_Q4;
assign R28C25_S27 = R28C25_Q7;
assign R28C25_N20 = R28C25_Q0;
assign R28C25_N23 = R28C25_Q3;
assign R28C25_S20 = R28C25_Q0;
assign R28C25_S23 = R28C25_Q3;
assign R28C25_N80 = R28C25_Q0;
assign R28C25_S80 = R28C25_Q0;
assign R28C25_E83 = R28C25_Q5;
assign R28C25_W83 = R28C25_Q5;
assign R28C25_E25 = R28C25_Q5;
assign R28C25_E26 = R28C25_Q6;
assign R28C25_W25 = R28C25_Q5;
assign R28C25_W26 = R28C25_Q6;
assign R28C25_E24 = R28C25_Q4;
assign R28C25_E27 = R28C25_Q7;
assign R28C25_W24 = R28C25_Q4;
assign R28C25_W27 = R28C25_Q7;
assign R28C25_E20 = R28C25_Q0;
assign R28C25_E23 = R28C25_Q3;
assign R28C25_W20 = R28C25_Q0;
assign R28C25_W23 = R28C25_Q3;
assign R28C25_B0 = R28C25_F3;
assign R28C25_B1 = R28C25_F3;
assign R28C25_B2 = R28C25_F1;
assign R28C25_B3 = R28C25_F1;
assign R28C25_B4 = R28C25_F1;
assign R28C25_B5 = R28C25_F1;
assign R28C25_B6 = R28C25_F1;
assign R28C25_B7 = R28C25_F1;
assign R28C25_D0 = R28C25_F2;
assign R28C25_D1 = R28C25_F2;
assign R28C25_D2 = R28C25_F0;
assign R28C25_D3 = R28C25_F0;
assign R28C25_D4 = R28C25_F0;
assign R28C25_D5 = R28C25_F0;
assign R28C25_D6 = R28C25_F0;
assign R28C25_D7 = R28C25_F0;
assign R28C25_X02 = R28C25_Q1;
assign R28C25_X04 = R28C25_Q7;
assign R28C25_X06 = R28C25_Q1;
assign R28C25_X08 = R28C25_Q7;
assign R28C25_X01 = R28C25_Q0;
assign R28C25_X03 = R28C25_Q6;
assign R28C25_X05 = R28C25_Q0;
assign R28C25_X07 = R28C25_Q6;
assign R28C25_N10 = R28C25_Q0;
assign R28C25_SN10 = R28C25_Q0;
assign R28C25_SN20 = R28C25_Q0;
assign R28C25_N13 = R28C25_Q0;
assign R28C25_S10 = R28C25_Q0;
assign R28C25_S13 = R28C25_Q0;
assign R28C25_E10 = R28C25_Q0;
assign R28C25_EW10 = R28C25_Q0;
assign R28C25_EW20 = R28C25_Q0;
assign R28C25_E13 = R28C25_Q0;
assign R28C25_W10 = R28C25_Q0;
assign R28C25_W13 = R28C25_Q0;
assign R28C25_E11 = R28C25_EW10;
assign R28C25_W11 = R28C25_EW10;
assign R28C25_E12 = R28C25_EW20;
assign R28C25_W12 = R28C25_EW20;
assign R28C25_S11 = R28C25_SN10;
assign R28C25_N11 = R28C25_SN10;
assign R28C25_S12 = R28C25_SN20;
assign R28C25_N12 = R28C25_SN20;
assign R28C28_CLK0 = VCC;
assign R28C28_CLK1 = VCC;
assign R28C28_CLK2 = VCC;
assign R28C28_LSR0 = VCC;
assign R28C28_LSR1 = VCC;
assign R28C28_LSR2 = VCC;
assign R28C28_CE0 = VCC;
assign R28C28_CE1 = VCC;
assign R28C28_CE2 = VCC;
assign R28C28_SEL0 = VCC;
assign R28C28_SEL1 = VCC;
assign R28C28_SEL2 = VCC;
assign R28C28_SEL3 = VCC;
assign R28C28_SEL4 = VCC;
assign R28C28_SEL5 = VCC;
assign R28C28_SEL6 = VCC;
assign R28C28_SEL7 = VCC;
assign R28C28_C0 = R28C28_F4;
assign R28C28_C1 = R28C28_F4;
assign R28C28_C2 = R28C28_F4;
assign R28C28_C3 = R28C28_F4;
assign R28C28_A4 = R28C28_F7;
assign R28C28_A5 = R28C28_F7;
assign R28C28_A6 = R28C28_F5;
assign R28C28_A7 = R28C28_F5;
assign R28C28_N82 = R28C28_Q4;
assign R28C28_S82 = R28C28_Q4;
assign R28C28_E82 = R28C28_Q4;
assign R28C28_W82 = R28C28_Q4;
assign R28C28_A0 = R28C28_F5;
assign R28C28_A1 = R28C28_F5;
assign R28C28_A2 = R28C28_F5;
assign R28C28_A3 = R28C28_F5;
assign R28C28_C4 = R28C28_F6;
assign R28C28_C5 = R28C28_F6;
assign R28C28_C6 = R28C28_F4;
assign R28C28_C7 = R28C28_F4;
assign R28C28_N81 = R28C28_Q1;
assign R28C28_S81 = R28C28_Q1;
assign R28C28_E81 = R28C28_Q1;
assign R28C28_W81 = R28C28_Q1;
assign R28C28_N21 = R28C28_Q1;
assign R28C28_N22 = R28C28_Q2;
assign R28C28_S21 = R28C28_Q1;
assign R28C28_S22 = R28C28_Q2;
assign R28C28_E21 = R28C28_Q1;
assign R28C28_E22 = R28C28_Q2;
assign R28C28_W21 = R28C28_Q1;
assign R28C28_W22 = R28C28_Q2;
assign R28C28_E80 = R28C28_Q0;
assign R28C28_W80 = R28C28_Q0;
assign R28C28_N25 = R28C28_Q5;
assign R28C28_N26 = R28C28_Q6;
assign R28C28_S25 = R28C28_Q5;
assign R28C28_S26 = R28C28_Q6;
assign R28C28_N83 = R28C28_Q5;
assign R28C28_S83 = R28C28_Q5;
assign R28C28_N24 = R28C28_Q4;
assign R28C28_N27 = R28C28_Q7;
assign R28C28_S24 = R28C28_Q4;
assign R28C28_S27 = R28C28_Q7;
assign R28C28_N20 = R28C28_Q0;
assign R28C28_N23 = R28C28_Q3;
assign R28C28_S20 = R28C28_Q0;
assign R28C28_S23 = R28C28_Q3;
assign R28C28_N80 = R28C28_Q0;
assign R28C28_S80 = R28C28_Q0;
assign R28C28_E83 = R28C28_Q5;
assign R28C28_W83 = R28C28_Q5;
assign R28C28_E25 = R28C28_Q5;
assign R28C28_E26 = R28C28_Q6;
assign R28C28_W25 = R28C28_Q5;
assign R28C28_W26 = R28C28_Q6;
assign R28C28_E24 = R28C28_Q4;
assign R28C28_E27 = R28C28_Q7;
assign R28C28_W24 = R28C28_Q4;
assign R28C28_W27 = R28C28_Q7;
assign R28C28_E20 = R28C28_Q0;
assign R28C28_E23 = R28C28_Q3;
assign R28C28_W20 = R28C28_Q0;
assign R28C28_W23 = R28C28_Q3;
assign R28C28_B0 = R28C28_F3;
assign R28C28_B1 = R28C28_F3;
assign R28C28_B2 = R28C28_F1;
assign R28C28_B3 = R28C28_F1;
assign R28C28_B4 = R28C28_F1;
assign R28C28_B5 = R28C28_F1;
assign R28C28_B6 = R28C28_F1;
assign R28C28_B7 = R28C28_F1;
assign R28C28_D0 = R28C28_F2;
assign R28C28_D1 = R28C28_F2;
assign R28C28_D2 = R28C28_F0;
assign R28C28_D3 = R28C28_F0;
assign R28C28_D4 = R28C28_F0;
assign R28C28_D5 = R28C28_F0;
assign R28C28_D6 = R28C28_F0;
assign R28C28_D7 = R28C28_F0;
assign R28C28_X02 = R28C28_Q1;
assign R28C28_X04 = R28C28_Q7;
assign R28C28_X06 = R28C28_Q1;
assign R28C28_X08 = R28C28_Q7;
assign R28C28_X01 = R28C28_Q0;
assign R28C28_X03 = R28C28_Q6;
assign R28C28_X05 = R28C28_Q0;
assign R28C28_X07 = R28C28_Q6;
assign R28C28_N10 = R28C28_Q0;
assign R28C28_SN10 = R28C28_Q0;
assign R28C28_SN20 = R28C28_Q0;
assign R28C28_N13 = R28C28_Q0;
assign R28C28_S10 = R28C28_Q0;
assign R28C28_S13 = R28C28_Q0;
assign R28C28_E10 = R28C28_Q0;
assign R28C28_EW10 = R28C28_Q0;
assign R28C28_EW20 = R28C28_Q0;
assign R28C28_E13 = R28C28_Q0;
assign R28C28_W10 = R28C28_Q0;
assign R28C28_W13 = R28C28_Q0;
assign R28C28_E11 = R28C28_EW10;
assign R28C28_W11 = R28C28_EW10;
assign R28C28_E12 = R28C28_EW20;
assign R28C28_W12 = R28C28_EW20;
assign R28C28_S11 = R28C28_SN10;
assign R28C28_N11 = R28C28_SN10;
assign R28C28_S12 = R28C28_SN20;
assign R28C28_N12 = R28C28_SN20;
assign R28C31_CLK0 = VCC;
assign R28C31_CLK1 = VCC;
assign R28C31_CLK2 = VCC;
assign R28C31_LSR0 = VCC;
assign R28C31_LSR1 = VCC;
assign R28C31_LSR2 = VCC;
assign R28C31_CE0 = VCC;
assign R28C31_CE1 = VCC;
assign R28C31_CE2 = VCC;
assign R28C31_SEL0 = VCC;
assign R28C31_SEL1 = VCC;
assign R28C31_SEL2 = VCC;
assign R28C31_SEL3 = VCC;
assign R28C31_SEL4 = VCC;
assign R28C31_SEL5 = VCC;
assign R28C31_SEL6 = VCC;
assign R28C31_SEL7 = VCC;
assign R28C31_C0 = R28C31_F4;
assign R28C31_C1 = R28C31_F4;
assign R28C31_C2 = R28C31_F4;
assign R28C31_C3 = R28C31_F4;
assign R28C31_A4 = R28C31_F7;
assign R28C31_A5 = R28C31_F7;
assign R28C31_A6 = R28C31_F5;
assign R28C31_A7 = R28C31_F5;
assign R28C31_N82 = R28C31_Q4;
assign R28C31_S82 = R28C31_Q4;
assign R28C31_E82 = R28C31_Q4;
assign R28C31_W82 = R28C31_Q4;
assign R28C31_A0 = R28C31_F5;
assign R28C31_A1 = R28C31_F5;
assign R28C31_A2 = R28C31_F5;
assign R28C31_A3 = R28C31_F5;
assign R28C31_C4 = R28C31_F6;
assign R28C31_C5 = R28C31_F6;
assign R28C31_C6 = R28C31_F4;
assign R28C31_C7 = R28C31_F4;
assign R28C31_N81 = R28C31_Q1;
assign R28C31_S81 = R28C31_Q1;
assign R28C31_E81 = R28C31_Q1;
assign R28C31_W81 = R28C31_Q1;
assign R28C31_N21 = R28C31_Q1;
assign R28C31_N22 = R28C31_Q2;
assign R28C31_S21 = R28C31_Q1;
assign R28C31_S22 = R28C31_Q2;
assign R28C31_E21 = R28C31_Q1;
assign R28C31_E22 = R28C31_Q2;
assign R28C31_W21 = R28C31_Q1;
assign R28C31_W22 = R28C31_Q2;
assign R28C31_E80 = R28C31_Q0;
assign R28C31_W80 = R28C31_Q0;
assign R28C31_N25 = R28C31_Q5;
assign R28C31_N26 = R28C31_Q6;
assign R28C31_S25 = R28C31_Q5;
assign R28C31_S26 = R28C31_Q6;
assign R28C31_N83 = R28C31_Q5;
assign R28C31_S83 = R28C31_Q5;
assign R28C31_N24 = R28C31_Q4;
assign R28C31_N27 = R28C31_Q7;
assign R28C31_S24 = R28C31_Q4;
assign R28C31_S27 = R28C31_Q7;
assign R28C31_N20 = R28C31_Q0;
assign R28C31_N23 = R28C31_Q3;
assign R28C31_S20 = R28C31_Q0;
assign R28C31_S23 = R28C31_Q3;
assign R28C31_N80 = R28C31_Q0;
assign R28C31_S80 = R28C31_Q0;
assign R28C31_E83 = R28C31_Q5;
assign R28C31_W83 = R28C31_Q5;
assign R28C31_E25 = R28C31_Q5;
assign R28C31_E26 = R28C31_Q6;
assign R28C31_W25 = R28C31_Q5;
assign R28C31_W26 = R28C31_Q6;
assign R28C31_E24 = R28C31_Q4;
assign R28C31_E27 = R28C31_Q7;
assign R28C31_W24 = R28C31_Q4;
assign R28C31_W27 = R28C31_Q7;
assign R28C31_E20 = R28C31_Q0;
assign R28C31_E23 = R28C31_Q3;
assign R28C31_W20 = R28C31_Q0;
assign R28C31_W23 = R28C31_Q3;
assign R28C31_B0 = R28C31_F3;
assign R28C31_B1 = R28C31_F3;
assign R28C31_B2 = R28C31_F1;
assign R28C31_B3 = R28C31_F1;
assign R28C31_B4 = R28C31_F1;
assign R28C31_B5 = R28C31_F1;
assign R28C31_B6 = R28C31_F1;
assign R28C31_B7 = R28C31_F1;
assign R28C31_D0 = R28C31_F2;
assign R28C31_D1 = R28C31_F2;
assign R28C31_D2 = R28C31_F0;
assign R28C31_D3 = R28C31_F0;
assign R28C31_D4 = R28C31_F0;
assign R28C31_D5 = R28C31_F0;
assign R28C31_D6 = R28C31_F0;
assign R28C31_D7 = R28C31_F0;
assign R28C31_X02 = R28C31_Q1;
assign R28C31_X04 = R28C31_Q7;
assign R28C31_X06 = R28C31_Q1;
assign R28C31_X08 = R28C31_Q7;
assign R28C31_X01 = R28C31_Q0;
assign R28C31_X03 = R28C31_Q6;
assign R28C31_X05 = R28C31_Q0;
assign R28C31_X07 = R28C31_Q6;
assign R28C31_N10 = R28C31_Q0;
assign R28C31_SN10 = R28C31_Q0;
assign R28C31_SN20 = R28C31_Q0;
assign R28C31_N13 = R28C31_Q0;
assign R28C31_S10 = R28C31_Q0;
assign R28C31_S13 = R28C31_Q0;
assign R28C31_E10 = R28C31_Q0;
assign R28C31_EW10 = R28C31_Q0;
assign R28C31_EW20 = R28C31_Q0;
assign R28C31_E13 = R28C31_Q0;
assign R28C31_W10 = R28C31_Q0;
assign R28C31_W13 = R28C31_Q0;
assign R28C31_E11 = R28C31_EW10;
assign R28C31_W11 = R28C31_EW10;
assign R28C31_E12 = R28C31_EW20;
assign R28C31_W12 = R28C31_EW20;
assign R28C31_S11 = R28C31_SN10;
assign R28C31_N11 = R28C31_SN10;
assign R28C31_S12 = R28C31_SN20;
assign R28C31_N12 = R28C31_SN20;
assign R28C34_CLK0 = VCC;
assign R28C34_CLK1 = VCC;
assign R28C34_CLK2 = VCC;
assign R28C34_LSR0 = VCC;
assign R28C34_LSR1 = VCC;
assign R28C34_LSR2 = VCC;
assign R28C34_CE0 = VCC;
assign R28C34_CE1 = VCC;
assign R28C34_CE2 = VCC;
assign R28C34_SEL0 = VCC;
assign R28C34_SEL1 = VCC;
assign R28C34_SEL2 = VCC;
assign R28C34_SEL3 = VCC;
assign R28C34_SEL4 = VCC;
assign R28C34_SEL5 = VCC;
assign R28C34_SEL6 = VCC;
assign R28C34_SEL7 = VCC;
assign R28C34_C0 = R28C34_F4;
assign R28C34_C1 = R28C34_F4;
assign R28C34_C2 = R28C34_F4;
assign R28C34_C3 = R28C34_F4;
assign R28C34_A4 = R28C34_F7;
assign R28C34_A5 = R28C34_F7;
assign R28C34_A6 = R28C34_F5;
assign R28C34_A7 = R28C34_F5;
assign R28C34_N82 = R28C34_Q4;
assign R28C34_S82 = R28C34_Q4;
assign R28C34_E82 = R28C34_Q4;
assign R28C34_W82 = R28C34_Q4;
assign R28C34_A0 = R28C34_F5;
assign R28C34_A1 = R28C34_F5;
assign R28C34_A2 = R28C34_F5;
assign R28C34_A3 = R28C34_F5;
assign R28C34_C4 = R28C34_F6;
assign R28C34_C5 = R28C34_F6;
assign R28C34_C6 = R28C34_F4;
assign R28C34_C7 = R28C34_F4;
assign R28C34_N81 = R28C34_Q1;
assign R28C34_S81 = R28C34_Q1;
assign R28C34_E81 = R28C34_Q1;
assign R28C34_W81 = R28C34_Q1;
assign R28C34_N21 = R28C34_Q1;
assign R28C34_N22 = R28C34_Q2;
assign R28C34_S21 = R28C34_Q1;
assign R28C34_S22 = R28C34_Q2;
assign R28C34_E21 = R28C34_Q1;
assign R28C34_E22 = R28C34_Q2;
assign R28C34_W21 = R28C34_Q1;
assign R28C34_W22 = R28C34_Q2;
assign R28C34_E80 = R28C34_Q0;
assign R28C34_W80 = R28C34_Q0;
assign R28C34_N25 = R28C34_Q5;
assign R28C34_N26 = R28C34_Q6;
assign R28C34_S25 = R28C34_Q5;
assign R28C34_S26 = R28C34_Q6;
assign R28C34_N83 = R28C34_Q5;
assign R28C34_S83 = R28C34_Q5;
assign R28C34_N24 = R28C34_Q4;
assign R28C34_N27 = R28C34_Q7;
assign R28C34_S24 = R28C34_Q4;
assign R28C34_S27 = R28C34_Q7;
assign R28C34_N20 = R28C34_Q0;
assign R28C34_N23 = R28C34_Q3;
assign R28C34_S20 = R28C34_Q0;
assign R28C34_S23 = R28C34_Q3;
assign R28C34_N80 = R28C34_Q0;
assign R28C34_S80 = R28C34_Q0;
assign R28C34_E83 = R28C34_Q5;
assign R28C34_W83 = R28C34_Q5;
assign R28C34_E25 = R28C34_Q5;
assign R28C34_E26 = R28C34_Q6;
assign R28C34_W25 = R28C34_Q5;
assign R28C34_W26 = R28C34_Q6;
assign R28C34_E24 = R28C34_Q4;
assign R28C34_E27 = R28C34_Q7;
assign R28C34_W24 = R28C34_Q4;
assign R28C34_W27 = R28C34_Q7;
assign R28C34_E20 = R28C34_Q0;
assign R28C34_E23 = R28C34_Q3;
assign R28C34_W20 = R28C34_Q0;
assign R28C34_W23 = R28C34_Q3;
assign R28C34_B0 = R28C34_F3;
assign R28C34_B1 = R28C34_F3;
assign R28C34_B2 = R28C34_F1;
assign R28C34_B3 = R28C34_F1;
assign R28C34_B4 = R28C34_F1;
assign R28C34_B5 = R28C34_F1;
assign R28C34_B6 = R28C34_F1;
assign R28C34_B7 = R28C34_F1;
assign R28C34_D0 = R28C34_F2;
assign R28C34_D1 = R28C34_F2;
assign R28C34_D2 = R28C34_F0;
assign R28C34_D3 = R28C34_F0;
assign R28C34_D4 = R28C34_F0;
assign R28C34_D5 = R28C34_F0;
assign R28C34_D6 = R28C34_F0;
assign R28C34_D7 = R28C34_F0;
assign R28C34_X02 = R28C34_Q1;
assign R28C34_X04 = R28C34_Q7;
assign R28C34_X06 = R28C34_Q1;
assign R28C34_X08 = R28C34_Q7;
assign R28C34_X01 = R28C34_Q0;
assign R28C34_X03 = R28C34_Q6;
assign R28C34_X05 = R28C34_Q0;
assign R28C34_X07 = R28C34_Q6;
assign R28C34_N10 = R28C34_Q0;
assign R28C34_SN10 = R28C34_Q0;
assign R28C34_SN20 = R28C34_Q0;
assign R28C34_N13 = R28C34_Q0;
assign R28C34_S10 = R28C34_Q0;
assign R28C34_S13 = R28C34_Q0;
assign R28C34_E10 = R28C34_Q0;
assign R28C34_EW10 = R28C34_Q0;
assign R28C34_EW20 = R28C34_Q0;
assign R28C34_E13 = R28C34_Q0;
assign R28C34_W10 = R28C34_Q0;
assign R28C34_W13 = R28C34_Q0;
assign R28C34_E11 = R28C34_EW10;
assign R28C34_W11 = R28C34_EW10;
assign R28C34_E12 = R28C34_EW20;
assign R28C34_W12 = R28C34_EW20;
assign R28C34_S11 = R28C34_SN10;
assign R28C34_N11 = R28C34_SN10;
assign R28C34_S12 = R28C34_SN20;
assign R28C34_N12 = R28C34_SN20;
assign R28C37_CLK0 = VCC;
assign R28C37_CLK1 = VCC;
assign R28C37_CLK2 = VCC;
assign R28C37_LSR0 = VCC;
assign R28C37_LSR1 = VCC;
assign R28C37_LSR2 = VCC;
assign R28C37_CE0 = VCC;
assign R28C37_CE1 = VCC;
assign R28C37_CE2 = VCC;
assign R28C37_SEL0 = VCC;
assign R28C37_SEL1 = VCC;
assign R28C37_SEL2 = VCC;
assign R28C37_SEL3 = VCC;
assign R28C37_SEL4 = VCC;
assign R28C37_SEL5 = VCC;
assign R28C37_SEL6 = VCC;
assign R28C37_SEL7 = VCC;
assign R28C37_C0 = R28C37_F4;
assign R28C37_C1 = R28C37_F4;
assign R28C37_C2 = R28C37_F4;
assign R28C37_C3 = R28C37_F4;
assign R28C37_A4 = R28C37_F7;
assign R28C37_A5 = R28C37_F7;
assign R28C37_A6 = R28C37_F5;
assign R28C37_A7 = R28C37_F5;
assign R28C37_N82 = R28C37_Q4;
assign R28C37_S82 = R28C37_Q4;
assign R28C37_E82 = R28C37_Q4;
assign R28C37_W82 = R28C37_Q4;
assign R28C37_A0 = R28C37_F5;
assign R28C37_A1 = R28C37_F5;
assign R28C37_A2 = R28C37_F5;
assign R28C37_A3 = R28C37_F5;
assign R28C37_C4 = R28C37_F6;
assign R28C37_C5 = R28C37_F6;
assign R28C37_C6 = R28C37_F4;
assign R28C37_C7 = R28C37_F4;
assign R28C37_N81 = R28C37_Q1;
assign R28C37_S81 = R28C37_Q1;
assign R28C37_E81 = R28C37_Q1;
assign R28C37_W81 = R28C37_Q1;
assign R28C37_N21 = R28C37_Q1;
assign R28C37_N22 = R28C37_Q2;
assign R28C37_S21 = R28C37_Q1;
assign R28C37_S22 = R28C37_Q2;
assign R28C37_E21 = R28C37_Q1;
assign R28C37_E22 = R28C37_Q2;
assign R28C37_W21 = R28C37_Q1;
assign R28C37_W22 = R28C37_Q2;
assign R28C37_E80 = R28C37_Q0;
assign R28C37_W80 = R28C37_Q0;
assign R28C37_N25 = R28C37_Q5;
assign R28C37_N26 = R28C37_Q6;
assign R28C37_S25 = R28C37_Q5;
assign R28C37_S26 = R28C37_Q6;
assign R28C37_N83 = R28C37_Q5;
assign R28C37_S83 = R28C37_Q5;
assign R28C37_N24 = R28C37_Q4;
assign R28C37_N27 = R28C37_Q7;
assign R28C37_S24 = R28C37_Q4;
assign R28C37_S27 = R28C37_Q7;
assign R28C37_N20 = R28C37_Q0;
assign R28C37_N23 = R28C37_Q3;
assign R28C37_S20 = R28C37_Q0;
assign R28C37_S23 = R28C37_Q3;
assign R28C37_N80 = R28C37_Q0;
assign R28C37_S80 = R28C37_Q0;
assign R28C37_E83 = R28C37_Q5;
assign R28C37_W83 = R28C37_Q5;
assign R28C37_E25 = R28C37_Q5;
assign R28C37_E26 = R28C37_Q6;
assign R28C37_W25 = R28C37_Q5;
assign R28C37_W26 = R28C37_Q6;
assign R28C37_E24 = R28C37_Q4;
assign R28C37_E27 = R28C37_Q7;
assign R28C37_W24 = R28C37_Q4;
assign R28C37_W27 = R28C37_Q7;
assign R28C37_E20 = R28C37_Q0;
assign R28C37_E23 = R28C37_Q3;
assign R28C37_W20 = R28C37_Q0;
assign R28C37_W23 = R28C37_Q3;
assign R28C37_B0 = R28C37_F3;
assign R28C37_B1 = R28C37_F3;
assign R28C37_B2 = R28C37_F1;
assign R28C37_B3 = R28C37_F1;
assign R28C37_B4 = R28C37_F1;
assign R28C37_B5 = R28C37_F1;
assign R28C37_B6 = R28C37_F1;
assign R28C37_B7 = R28C37_F1;
assign R28C37_D0 = R28C37_F2;
assign R28C37_D1 = R28C37_F2;
assign R28C37_D2 = R28C37_F0;
assign R28C37_D3 = R28C37_F0;
assign R28C37_D4 = R28C37_F0;
assign R28C37_D5 = R28C37_F0;
assign R28C37_D6 = R28C37_F0;
assign R28C37_D7 = R28C37_F0;
assign R28C37_X02 = R28C37_Q1;
assign R28C37_X04 = R28C37_Q7;
assign R28C37_X06 = R28C37_Q1;
assign R28C37_X08 = R28C37_Q7;
assign R28C37_X01 = R28C37_Q0;
assign R28C37_X03 = R28C37_Q6;
assign R28C37_X05 = R28C37_Q0;
assign R28C37_X07 = R28C37_Q6;
assign R28C37_N10 = R28C37_Q0;
assign R28C37_SN10 = R28C37_Q0;
assign R28C37_SN20 = R28C37_Q0;
assign R28C37_N13 = R28C37_Q0;
assign R28C37_S10 = R28C37_Q0;
assign R28C37_S13 = R28C37_Q0;
assign R28C37_E10 = R28C37_Q0;
assign R28C37_EW10 = R28C37_Q0;
assign R28C37_EW20 = R28C37_Q0;
assign R28C37_E13 = R28C37_Q0;
assign R28C37_W10 = R28C37_Q0;
assign R28C37_W13 = R28C37_Q0;
assign R28C37_E11 = R28C37_EW10;
assign R28C37_W11 = R28C37_EW10;
assign R28C37_E12 = R28C37_EW20;
assign R28C37_W12 = R28C37_EW20;
assign R28C37_S11 = R28C37_SN10;
assign R28C37_N11 = R28C37_SN10;
assign R28C37_S12 = R28C37_SN20;
assign R28C37_N12 = R28C37_SN20;
assign R28C40_CLK0 = VCC;
assign R28C40_CLK1 = VCC;
assign R28C40_CLK2 = VCC;
assign R28C40_LSR0 = VCC;
assign R28C40_LSR1 = VCC;
assign R28C40_LSR2 = VCC;
assign R28C40_CE0 = VCC;
assign R28C40_CE1 = VCC;
assign R28C40_CE2 = VCC;
assign R28C40_SEL0 = VCC;
assign R28C40_SEL1 = VCC;
assign R28C40_SEL2 = VCC;
assign R28C40_SEL3 = VCC;
assign R28C40_SEL4 = VCC;
assign R28C40_SEL5 = VCC;
assign R28C40_SEL6 = VCC;
assign R28C40_SEL7 = VCC;
assign R28C40_C0 = R28C40_F4;
assign R28C40_C1 = R28C40_F4;
assign R28C40_C2 = R28C40_F4;
assign R28C40_C3 = R28C40_F4;
assign R28C40_A4 = R28C40_F7;
assign R28C40_A5 = R28C40_F7;
assign R28C40_A6 = R28C40_F5;
assign R28C40_A7 = R28C40_F5;
assign R28C40_N82 = R28C40_Q4;
assign R28C40_S82 = R28C40_Q4;
assign R28C40_E82 = R28C40_Q4;
assign R28C40_W82 = R28C40_Q4;
assign R28C40_A0 = R28C40_F5;
assign R28C40_A1 = R28C40_F5;
assign R28C40_A2 = R28C40_F5;
assign R28C40_A3 = R28C40_F5;
assign R28C40_C4 = R28C40_F6;
assign R28C40_C5 = R28C40_F6;
assign R28C40_C6 = R28C40_F4;
assign R28C40_C7 = R28C40_F4;
assign R28C40_N81 = R28C40_Q1;
assign R28C40_S81 = R28C40_Q1;
assign R28C40_E81 = R28C40_Q1;
assign R28C40_W81 = R28C40_Q1;
assign R28C40_N21 = R28C40_Q1;
assign R28C40_N22 = R28C40_Q2;
assign R28C40_S21 = R28C40_Q1;
assign R28C40_S22 = R28C40_Q2;
assign R28C40_E21 = R28C40_Q1;
assign R28C40_E22 = R28C40_Q2;
assign R28C40_W21 = R28C40_Q1;
assign R28C40_W22 = R28C40_Q2;
assign R28C40_E80 = R28C40_Q0;
assign R28C40_W80 = R28C40_Q0;
assign R28C40_N25 = R28C40_Q5;
assign R28C40_N26 = R28C40_Q6;
assign R28C40_S25 = R28C40_Q5;
assign R28C40_S26 = R28C40_Q6;
assign R28C40_N83 = R28C40_Q5;
assign R28C40_S83 = R28C40_Q5;
assign R28C40_N24 = R28C40_Q4;
assign R28C40_N27 = R28C40_Q7;
assign R28C40_S24 = R28C40_Q4;
assign R28C40_S27 = R28C40_Q7;
assign R28C40_N20 = R28C40_Q0;
assign R28C40_N23 = R28C40_Q3;
assign R28C40_S20 = R28C40_Q0;
assign R28C40_S23 = R28C40_Q3;
assign R28C40_N80 = R28C40_Q0;
assign R28C40_S80 = R28C40_Q0;
assign R28C40_E83 = R28C40_Q5;
assign R28C40_W83 = R28C40_Q5;
assign R28C40_E25 = R28C40_Q5;
assign R28C40_E26 = R28C40_Q6;
assign R28C40_W25 = R28C40_Q5;
assign R28C40_W26 = R28C40_Q6;
assign R28C40_E24 = R28C40_Q4;
assign R28C40_E27 = R28C40_Q7;
assign R28C40_W24 = R28C40_Q4;
assign R28C40_W27 = R28C40_Q7;
assign R28C40_E20 = R28C40_Q0;
assign R28C40_E23 = R28C40_Q3;
assign R28C40_W20 = R28C40_Q0;
assign R28C40_W23 = R28C40_Q3;
assign R28C40_B0 = R28C40_F3;
assign R28C40_B1 = R28C40_F3;
assign R28C40_B2 = R28C40_F1;
assign R28C40_B3 = R28C40_F1;
assign R28C40_B4 = R28C40_F1;
assign R28C40_B5 = R28C40_F1;
assign R28C40_B6 = R28C40_F1;
assign R28C40_B7 = R28C40_F1;
assign R28C40_D0 = R28C40_F2;
assign R28C40_D1 = R28C40_F2;
assign R28C40_D2 = R28C40_F0;
assign R28C40_D3 = R28C40_F0;
assign R28C40_D4 = R28C40_F0;
assign R28C40_D5 = R28C40_F0;
assign R28C40_D6 = R28C40_F0;
assign R28C40_D7 = R28C40_F0;
assign R28C40_X02 = R28C40_Q1;
assign R28C40_X04 = R28C40_Q7;
assign R28C40_X06 = R28C40_Q1;
assign R28C40_X08 = R28C40_Q7;
assign R28C40_X01 = R28C40_Q0;
assign R28C40_X03 = R28C40_Q6;
assign R28C40_X05 = R28C40_Q0;
assign R28C40_X07 = R28C40_Q6;
assign R28C40_N10 = R28C40_Q0;
assign R28C40_SN10 = R28C40_Q0;
assign R28C40_SN20 = R28C40_Q0;
assign R28C40_N13 = R28C40_Q0;
assign R28C40_S10 = R28C40_Q0;
assign R28C40_S13 = R28C40_Q0;
assign R28C40_E10 = R28C40_Q0;
assign R28C40_EW10 = R28C40_Q0;
assign R28C40_EW20 = R28C40_Q0;
assign R28C40_E13 = R28C40_Q0;
assign R28C40_W10 = R28C40_Q0;
assign R28C40_W13 = R28C40_Q0;
assign R28C40_E11 = R28C40_EW10;
assign R28C40_W11 = R28C40_EW10;
assign R28C40_E12 = R28C40_EW20;
assign R28C40_W12 = R28C40_EW20;
assign R28C40_S11 = R28C40_SN10;
assign R28C40_N11 = R28C40_SN10;
assign R28C40_S12 = R28C40_SN20;
assign R28C40_N12 = R28C40_SN20;
assign R28C43_CLK0 = VCC;
assign R28C43_CLK1 = VCC;
assign R28C43_CLK2 = VCC;
assign R28C43_LSR0 = VCC;
assign R28C43_LSR1 = VCC;
assign R28C43_LSR2 = VCC;
assign R28C43_CE0 = VCC;
assign R28C43_CE1 = VCC;
assign R28C43_CE2 = VCC;
assign R28C43_SEL0 = VCC;
assign R28C43_SEL1 = VCC;
assign R28C43_SEL2 = VCC;
assign R28C43_SEL3 = VCC;
assign R28C43_SEL4 = VCC;
assign R28C43_SEL5 = VCC;
assign R28C43_SEL6 = VCC;
assign R28C43_SEL7 = VCC;
assign R28C43_C0 = R28C43_F4;
assign R28C43_C1 = R28C43_F4;
assign R28C43_C2 = R28C43_F4;
assign R28C43_C3 = R28C43_F4;
assign R28C43_A4 = R28C43_F7;
assign R28C43_A5 = R28C43_F7;
assign R28C43_A6 = R28C43_F5;
assign R28C43_A7 = R28C43_F5;
assign R28C43_N82 = R28C43_Q4;
assign R28C43_S82 = R28C43_Q4;
assign R28C43_E82 = R28C43_Q4;
assign R28C43_W82 = R28C43_Q4;
assign R28C43_A0 = R28C43_F5;
assign R28C43_A1 = R28C43_F5;
assign R28C43_A2 = R28C43_F5;
assign R28C43_A3 = R28C43_F5;
assign R28C43_C4 = R28C43_F6;
assign R28C43_C5 = R28C43_F6;
assign R28C43_C6 = R28C43_F4;
assign R28C43_C7 = R28C43_F4;
assign R28C43_N81 = R28C43_Q1;
assign R28C43_S81 = R28C43_Q1;
assign R28C43_E81 = R28C43_Q1;
assign R28C43_W81 = R28C43_Q1;
assign R28C43_N21 = R28C43_Q1;
assign R28C43_N22 = R28C43_Q2;
assign R28C43_S21 = R28C43_Q1;
assign R28C43_S22 = R28C43_Q2;
assign R28C43_E21 = R28C43_Q1;
assign R28C43_E22 = R28C43_Q2;
assign R28C43_W21 = R28C43_Q1;
assign R28C43_W22 = R28C43_Q2;
assign R28C43_E80 = R28C43_Q0;
assign R28C43_W80 = R28C43_Q0;
assign R28C43_N25 = R28C43_Q5;
assign R28C43_N26 = R28C43_Q6;
assign R28C43_S25 = R28C43_Q5;
assign R28C43_S26 = R28C43_Q6;
assign R28C43_N83 = R28C43_Q5;
assign R28C43_S83 = R28C43_Q5;
assign R28C43_N24 = R28C43_Q4;
assign R28C43_N27 = R28C43_Q7;
assign R28C43_S24 = R28C43_Q4;
assign R28C43_S27 = R28C43_Q7;
assign R28C43_N20 = R28C43_Q0;
assign R28C43_N23 = R28C43_Q3;
assign R28C43_S20 = R28C43_Q0;
assign R28C43_S23 = R28C43_Q3;
assign R28C43_N80 = R28C43_Q0;
assign R28C43_S80 = R28C43_Q0;
assign R28C43_E83 = R28C43_Q5;
assign R28C43_W83 = R28C43_Q5;
assign R28C43_E25 = R28C43_Q5;
assign R28C43_E26 = R28C43_Q6;
assign R28C43_W25 = R28C43_Q5;
assign R28C43_W26 = R28C43_Q6;
assign R28C43_E24 = R28C43_Q4;
assign R28C43_E27 = R28C43_Q7;
assign R28C43_W24 = R28C43_Q4;
assign R28C43_W27 = R28C43_Q7;
assign R28C43_E20 = R28C43_Q0;
assign R28C43_E23 = R28C43_Q3;
assign R28C43_W20 = R28C43_Q0;
assign R28C43_W23 = R28C43_Q3;
assign R28C43_B0 = R28C43_F3;
assign R28C43_B1 = R28C43_F3;
assign R28C43_B2 = R28C43_F1;
assign R28C43_B3 = R28C43_F1;
assign R28C43_B4 = R28C43_F1;
assign R28C43_B5 = R28C43_F1;
assign R28C43_B6 = R28C43_F1;
assign R28C43_B7 = R28C43_F1;
assign R28C43_D0 = R28C43_F2;
assign R28C43_D1 = R28C43_F2;
assign R28C43_D2 = R28C43_F0;
assign R28C43_D3 = R28C43_F0;
assign R28C43_D4 = R28C43_F0;
assign R28C43_D5 = R28C43_F0;
assign R28C43_D6 = R28C43_F0;
assign R28C43_D7 = R28C43_F0;
assign R28C43_X02 = R28C43_Q1;
assign R28C43_X04 = R28C43_Q7;
assign R28C43_X06 = R28C43_Q1;
assign R28C43_X08 = R28C43_Q7;
assign R28C43_X01 = R28C43_Q0;
assign R28C43_X03 = R28C43_Q6;
assign R28C43_X05 = R28C43_Q0;
assign R28C43_X07 = R28C43_Q6;
assign R28C43_N10 = R28C43_Q0;
assign R28C43_SN10 = R28C43_Q0;
assign R28C43_SN20 = R28C43_Q0;
assign R28C43_N13 = R28C43_Q0;
assign R28C43_S10 = R28C43_Q0;
assign R28C43_S13 = R28C43_Q0;
assign R28C43_E10 = R28C43_Q0;
assign R28C43_EW10 = R28C43_Q0;
assign R28C43_EW20 = R28C43_Q0;
assign R28C43_E13 = R28C43_Q0;
assign R28C43_W10 = R28C43_Q0;
assign R28C43_W13 = R28C43_Q0;
assign R28C43_E11 = R28C43_EW10;
assign R28C43_W11 = R28C43_EW10;
assign R28C43_E12 = R28C43_EW20;
assign R28C43_W12 = R28C43_EW20;
assign R28C43_S11 = R28C43_SN10;
assign R28C43_N11 = R28C43_SN10;
assign R28C43_S12 = R28C43_SN20;
assign R28C43_N12 = R28C43_SN20;
assign R28C46_CLK0 = VCC;
assign R28C46_CLK1 = VCC;
assign R28C46_CLK2 = VCC;
assign R28C46_LSR0 = VCC;
assign R28C46_LSR1 = VCC;
assign R28C46_LSR2 = VCC;
assign R28C46_CE0 = VCC;
assign R28C46_CE1 = VCC;
assign R28C46_CE2 = VCC;
assign R28C46_SEL0 = VCC;
assign R28C46_SEL1 = VCC;
assign R28C46_SEL2 = VCC;
assign R28C46_SEL3 = VCC;
assign R28C46_SEL4 = VCC;
assign R28C46_SEL5 = VCC;
assign R28C46_SEL6 = VCC;
assign R28C46_SEL7 = VCC;
assign R28C46_C0 = R28C46_F4;
assign R28C46_C1 = R28C46_F4;
assign R28C46_C2 = R28C46_F4;
assign R28C46_C3 = R28C46_F4;
assign R28C46_A4 = R28C46_F7;
assign R28C46_A5 = R28C46_F7;
assign R28C46_A6 = R28C46_F5;
assign R28C46_A7 = R28C46_F5;
assign R28C46_N82 = R28C46_Q4;
assign R28C46_S82 = R28C46_Q4;
assign R28C46_E82 = R28C46_Q4;
assign R28C46_W82 = R28C46_Q4;
assign R28C46_A0 = R28C46_F5;
assign R28C46_A1 = R28C46_F5;
assign R28C46_A2 = R28C46_F5;
assign R28C46_A3 = R28C46_F5;
assign R28C46_C4 = R28C46_F6;
assign R28C46_C5 = R28C46_F6;
assign R28C46_C6 = R28C46_F4;
assign R28C46_C7 = R28C46_F4;
assign R28C46_N81 = R28C46_Q1;
assign R28C46_S81 = R28C46_Q1;
assign R28C46_E81 = R28C46_Q1;
assign R28C46_W81 = R28C46_Q1;
assign R28C46_N21 = R28C46_Q1;
assign R28C46_N22 = R28C46_Q2;
assign R28C46_S21 = R28C46_Q1;
assign R28C46_S22 = R28C46_Q2;
assign R28C46_E21 = R28C46_Q1;
assign R28C46_E22 = R28C46_Q2;
assign R28C46_W21 = R28C46_Q1;
assign R28C46_W22 = R28C46_Q2;
assign R28C46_E80 = R28C46_Q0;
assign R28C46_W80 = R28C46_Q0;
assign R28C46_N25 = R28C46_Q5;
assign R28C46_N26 = R28C46_Q6;
assign R28C46_S25 = R28C46_Q5;
assign R28C46_S26 = R28C46_Q6;
assign R28C46_N83 = R28C46_Q5;
assign R28C46_S83 = R28C46_Q5;
assign R28C46_N24 = R28C46_Q4;
assign R28C46_N27 = R28C46_Q7;
assign R28C46_S24 = R28C46_Q4;
assign R28C46_S27 = R28C46_Q7;
assign R28C46_N20 = R28C46_Q0;
assign R28C46_N23 = R28C46_Q3;
assign R28C46_S20 = R28C46_Q0;
assign R28C46_S23 = R28C46_Q3;
assign R28C46_N80 = R28C46_Q0;
assign R28C46_S80 = R28C46_Q0;
assign R28C46_E83 = R28C46_Q5;
assign R28C46_W83 = R28C46_Q5;
assign R28C46_E25 = R28C46_Q5;
assign R28C46_E26 = R28C46_Q6;
assign R28C46_W25 = R28C46_Q5;
assign R28C46_W26 = R28C46_Q6;
assign R28C46_E24 = R28C46_Q4;
assign R28C46_E27 = R28C46_Q7;
assign R28C46_W24 = R28C46_Q4;
assign R28C46_W27 = R28C46_Q7;
assign R28C46_E20 = R28C46_Q0;
assign R28C46_E23 = R28C46_Q3;
assign R28C46_W20 = R28C46_Q0;
assign R28C46_W23 = R28C46_Q3;
assign R28C46_B0 = R28C46_F3;
assign R28C46_B1 = R28C46_F3;
assign R28C46_B2 = R28C46_F1;
assign R28C46_B3 = R28C46_F1;
assign R28C46_B4 = R28C46_F1;
assign R28C46_B5 = R28C46_F1;
assign R28C46_B6 = R28C46_F1;
assign R28C46_B7 = R28C46_F1;
assign R28C46_D0 = R28C46_F2;
assign R28C46_D1 = R28C46_F2;
assign R28C46_D2 = R28C46_F0;
assign R28C46_D3 = R28C46_F0;
assign R28C46_D4 = R28C46_F0;
assign R28C46_D5 = R28C46_F0;
assign R28C46_D6 = R28C46_F0;
assign R28C46_D7 = R28C46_F0;
assign R28C46_X02 = R28C46_Q1;
assign R28C46_X04 = R28C46_Q7;
assign R28C46_X06 = R28C46_Q1;
assign R28C46_X08 = R28C46_Q7;
assign R28C46_X01 = R28C46_Q0;
assign R28C46_X03 = R28C46_Q6;
assign R28C46_X05 = R28C46_Q0;
assign R28C46_X07 = R28C46_Q6;
assign R28C46_N10 = R28C46_Q0;
assign R28C46_SN10 = R28C46_Q0;
assign R28C46_SN20 = R28C46_Q0;
assign R28C46_N13 = R28C46_Q0;
assign R28C46_S10 = R28C46_Q0;
assign R28C46_S13 = R28C46_Q0;
assign R28C46_E10 = R28C46_Q0;
assign R28C46_EW10 = R28C46_Q0;
assign R28C46_EW20 = R28C46_Q0;
assign R28C46_E13 = R28C46_Q0;
assign R28C46_W10 = R28C46_Q0;
assign R28C46_W13 = R28C46_Q0;
assign R28C46_E11 = R28C46_EW10;
assign R28C46_W11 = R28C46_EW10;
assign R28C46_E12 = R28C46_EW20;
assign R28C46_W12 = R28C46_EW20;
assign R28C46_S11 = R28C46_SN10;
assign R28C46_N11 = R28C46_SN10;
assign R28C46_S12 = R28C46_SN20;
assign R28C46_N12 = R28C46_SN20;
assign R29C28_CLK0 = VCC;
assign R29C28_CLK1 = VCC;
assign R29C28_CLK2 = VCC;
assign R29C28_LSR0 = VCC;
assign R29C28_LSR1 = VCC;
assign R29C28_LSR2 = VCC;
assign R29C28_CE0 = VCC;
assign R29C28_CE1 = VCC;
assign R29C28_CE2 = VCC;
assign R29C28_SEL0 = VCC;
assign R29C28_SEL1 = VCC;
assign R29C28_SEL2 = VCC;
assign R29C28_SEL3 = VCC;
assign R29C28_SEL4 = VCC;
assign R29C28_SEL5 = VCC;
assign R29C28_SEL6 = VCC;
assign R29C28_SEL7 = VCC;
assign R29C28_C0 = R29C28_F4;
assign R29C28_C1 = R29C28_F4;
assign R29C28_C2 = R29C28_F4;
assign R29C28_C3 = R29C28_F4;
assign R29C28_A4 = R29C28_F7;
assign R29C28_A5 = R29C28_F7;
assign R29C28_A6 = R29C28_F5;
assign R29C28_A7 = R29C28_F5;
assign R29C28_N82 = R29C28_Q4;
assign R29C28_S82 = R29C28_Q4;
assign R29C28_E82 = R29C28_Q4;
assign R29C28_W82 = R29C28_Q4;
assign R29C28_A0 = R29C28_F5;
assign R29C28_A1 = R29C28_F5;
assign R29C28_A2 = R29C28_F5;
assign R29C28_A3 = R29C28_F5;
assign R29C28_C4 = R29C28_F6;
assign R29C28_C5 = R29C28_F6;
assign R29C28_C6 = R29C28_F4;
assign R29C28_C7 = R29C28_F4;
assign R29C28_N81 = R29C28_Q1;
assign R29C28_S81 = R29C28_Q1;
assign R29C28_E81 = R29C28_Q1;
assign R29C28_W81 = R29C28_Q1;
assign R29C28_N21 = R29C28_Q1;
assign R29C28_N22 = R29C28_Q2;
assign R29C28_S21 = R29C28_Q1;
assign R29C28_S22 = R29C28_Q2;
assign R29C28_E21 = R29C28_Q1;
assign R29C28_E22 = R29C28_Q2;
assign R29C28_W21 = R29C28_Q1;
assign R29C28_W22 = R29C28_Q2;
assign R29C28_E80 = R29C28_Q0;
assign R29C28_W80 = R29C28_Q0;
assign R29C28_N25 = R29C28_Q5;
assign R29C28_N26 = R29C28_Q6;
assign R29C28_S25 = R29C28_Q5;
assign R29C28_S26 = R29C28_Q6;
assign R29C28_N83 = R29C28_Q5;
assign R29C28_S83 = R29C28_Q5;
assign R29C28_N24 = R29C28_Q4;
assign R29C28_N27 = R29C28_Q7;
assign R29C28_S24 = R29C28_Q4;
assign R29C28_S27 = R29C28_Q7;
assign R29C28_N20 = R29C28_Q0;
assign R29C28_N23 = R29C28_Q3;
assign R29C28_S20 = R29C28_Q0;
assign R29C28_S23 = R29C28_Q3;
assign R29C28_N80 = R29C28_Q0;
assign R29C28_S80 = R29C28_Q0;
assign R29C28_E83 = R29C28_Q5;
assign R29C28_W83 = R29C28_Q5;
assign R29C28_E25 = R29C28_Q5;
assign R29C28_E26 = R29C28_Q6;
assign R29C28_W25 = R29C28_Q5;
assign R29C28_W26 = R29C28_Q6;
assign R29C28_E24 = R29C28_Q4;
assign R29C28_E27 = R29C28_Q7;
assign R29C28_W24 = R29C28_Q4;
assign R29C28_W27 = R29C28_Q7;
assign R29C28_E20 = R29C28_Q0;
assign R29C28_E23 = R29C28_Q3;
assign R29C28_W20 = R29C28_Q0;
assign R29C28_W23 = R29C28_Q3;
assign R29C28_B0 = R29C28_F3;
assign R29C28_B1 = R29C28_F3;
assign R29C28_B2 = R29C28_F1;
assign R29C28_B3 = R29C28_F1;
assign R29C28_B4 = R29C28_F1;
assign R29C28_B5 = R29C28_F1;
assign R29C28_B6 = R29C28_F1;
assign R29C28_B7 = R29C28_F1;
assign R29C28_D0 = R29C28_F2;
assign R29C28_D1 = R29C28_F2;
assign R29C28_D2 = R29C28_F0;
assign R29C28_D3 = R29C28_F0;
assign R29C28_D4 = R29C28_F0;
assign R29C28_D5 = R29C28_F0;
assign R29C28_D6 = R29C28_F0;
assign R29C28_D7 = R29C28_F0;
assign R29C28_X02 = R29C28_Q1;
assign R29C28_X04 = R29C28_Q7;
assign R29C28_X06 = R29C28_Q1;
assign R29C28_X08 = R29C28_Q7;
assign R29C28_X01 = R29C28_Q0;
assign R29C28_X03 = R29C28_Q6;
assign R29C28_X05 = R29C28_Q0;
assign R29C28_X07 = R29C28_Q6;
assign R29C28_N10 = R29C28_Q0;
assign R29C28_SN10 = R29C28_Q0;
assign R29C28_SN20 = R29C28_Q0;
assign R29C28_N13 = R29C28_Q0;
assign R29C28_S10 = R29C28_Q0;
assign R29C28_S13 = R29C28_Q0;
assign R29C28_E10 = R29C28_Q0;
assign R29C28_EW10 = R29C28_Q0;
assign R29C28_EW20 = R29C28_Q0;
assign R29C28_E13 = R29C28_Q0;
assign R29C28_W10 = R29C28_Q0;
assign R29C28_W13 = R29C28_Q0;
assign R29C28_E11 = R29C28_EW10;
assign R29C28_W11 = R29C28_EW10;
assign R29C28_E12 = R29C28_EW20;
assign R29C28_W12 = R29C28_EW20;
assign R29C28_S11 = R29C28_SN10;
assign R29C28_N11 = R29C28_SN10;
assign R29C28_S12 = R29C28_SN20;
assign R29C28_N12 = R29C28_SN20;
IOBUF R1C32_IOBUF_A (
.O(R1C32_F6),
.OEN(R1C32_B0),
.I(R1C32_A0),
.IO(R1C32_IOA)
);
endmodule
