../img-video-ram.vh