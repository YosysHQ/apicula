`define PLL_DYN
`define PLL_DEVICE "GW1NZ-1"
`define PLL_FCLKIN "27"
`define PLL_ODIV_SEL  8

`define PLL_FBDIV_SEL 15
`define PLL_IDIV_SEL  7

`define PLL_FBDIV_SEL_1 23
`define PLL_IDIV_SEL_1  7

