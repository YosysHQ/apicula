`ifndef _img3_vh_
`define _img3_vh_
    defparam rom3.INIT_RAM_00 = 288'h000000000000008CD48C45A25128944A29168C452210C8644221148B462311C8E47A3D20;
    defparam rom3.INIT_RAM_01 = 288'h8542A150A85432190C86432190A8542A190C8845231148843221146A1180000000000000;
    defparam rom3.INIT_RAM_02 = 288'h000000000000000000223C229148A4522D188E462210C8643219108C472391C8E47A4926;
    defparam rom3.INIT_RAM_03 = 288'h8542A150C86432190C86432190C86432190C88462391888431D042000000000000000000;
    defparam rom3.INIT_RAM_04 = 288'h00000000000000000000081E1128944A29188E46229108844221148C472391C8E47A4926;
    defparam rom3.INIT_RAM_05 = 288'h8542A150C86432190C8743A1D10884421D0E894523114863A04000000000000000000000;
    defparam rom3.INIT_RAM_06 = 288'h6B359ADFEFF7FAFC7E0000040EC8743A25188E47231188C46231188F47A3D1C8E47A4926;
    defparam rom3.INIT_RAM_07 = 288'h8542A150C86432190E8844A29168C45A29128844A210C74080000C3D1E9ACD66B51A8D46;
    defparam rom3.INIT_RAM_08 = 288'h6B359ADFEFF7FBFDFEBF0F800207443221188E472391C8E472391C8F47A3D1C8E47A4926;
    defparam rom3.INIT_RAM_09 = 288'h8542A150C86432190E894522D188E4622D148943A18E810000186A3D1E9ACD66B51A8D46;
    defparam rom3.INIT_RAM_0A = 288'h6B3D3ADFEFF7FBFDFEFF6F87C00103A221188E47231188C462311A8F47A3D1A8C4723D20;
    defparam rom3.INIT_RAM_0B = 288'h86432150A8542A150C884522D188E4622D1489439D02000030D47A43329ACD66B51A6CE4;
    defparam rom3.INIT_RAM_0C = 288'h6B6BBFDFEFF7FBFDFEFF7FB7C3E00081E1188E4622910894522D188D47A35188B45A3118;
    defparam rom3.INIT_RAM_0D = 288'h8843A190A8542A150C430000000113D22D14893B0400000168F47A5F359AD28A3431ACD6;
    defparam rom3.INIT_RAM_0E = 288'h8B7FBFDFEFF7FBFDFEFF7FBFDFE00000451C8E462210C8744A29168D47A35168A4522914;
    defparam rom3.INIT_RAM_0F = 288'h8A442190A8542A150A00000000000081E1147808000000E1E8F4926B359E146A3359ACD6;
    defparam rom3.INIT_RAM_10 = 288'hD77FBFDFEFF7FBFDFEFF7FB7C3E0000001188C45A2910894522D188D47A35188B45A3118;
    defparam rom3.INIT_RAM_11 = 288'h8943A1D0C8642A150A0000000000000041141000000002D1E8F4BE6B35A5146A3359ACD6;
    defparam rom3.INIT_RAM_12 = 288'hFF7FBFDFEFF7FBFDFEFF6F87C000000001168B4622D188C46A31188E47239188C4723D20;
    defparam rom3.INIT_RAM_13 = 288'h874421D1087432150A0000000A28E09800000000000002D1E8F4D66B35A8D46A3359ACD6;
    defparam rom3.INIT_RAM_14 = 288'hFF7FBFDFEFF7FBFDFEFF00000000000001148A45A351E8F472391C8E472391C8E47A4926;
    defparam rom3.INIT_RAM_15 = 288'h8643A25148943A190C10000011CA347000000000000000E1E8F4D66B35A8D46A3359ACD6;
    defparam rom3.INIT_RAM_16 = 288'hFF7FBFDFEFF7FBFDFEFF6F87C000000001148A45A351E8F46A31188E47239188C4724524;
    defparam rom3.INIT_RAM_17 = 288'h8643A21128843A190C7408000268E51A382600000000000168F4A86B35A8D46A3359ACD6;
    defparam rom3.INIT_RAM_18 = 288'hD77FBFDFEFF7FBFDFEFF7FB7C3E0000001148A45A351E8D4622D188D47A35188B462391E;
    defparam rom3.INIT_RAM_19 = 288'h864321D0E87432190C8632000000028A8D1C13000000000030D47A3D1EA8D46A3359ACD6;
    defparam rom3.INIT_RAM_1A = 288'h8B7FBFDFEFF7FBFDFEFF7FBFDFE0000001148A45A351E8D45A29168D47A35168A45A311C;
    defparam rom3.INIT_RAM_1B = 288'h86432190C86432190C864308400000028D468E140000000000186A3D1EA8D46A3359ACD6;
    defparam rom3.INIT_RAM_1C = 288'h6B6BBFDFEFF7FBFDFEFF7FBFDFE0000001168B462351E8D4622D188C46A31188B462311C;
    defparam rom3.INIT_RAM_1D = 288'h8743A1D0E8742A150A864319000000028D469B4998C4000000000C3D1EA8D469B389C4D6;
    defparam rom3.INIT_RAM_1E = 288'h6B3D3ADFEFF7FBFDFEFF772150A2000000D48D46A3D1E8F46A35188C45A31188C462391C;
    defparam rom3.INIT_RAM_1F = 288'h8944A251287432150A854321800000028D469B462150A631000000000028D469B429F8F0;
    defparam rom3.INIT_RAM_20 = 288'h71359E9AEFF7FBFDFEDD48A150A6300000468F47A3D1E8F47A3D1A8B4522D188E472391C;
    defparam rom3.INIT_RAM_21 = 288'h8A452291488432150A854321800000028D469B462150A854298C200009A8D469B46214FC;
    defparam rom3.INIT_RAM_22 = 288'h78389C4F09F6EB753E85429F9189314000006B47A3D1E8F46A35188B4522D188C462391C;
    defparam rom3.INIT_RAM_23 = 288'h8944A25128742A150A854310800000026D369349A31188C46214E61024A6D469B49A310A;
    defparam rom3.INIT_RAM_24 = 288'h853F1F8FC8542A150A853C1C4E29B4704C002347A3D1E8D4622D168A45229168B462311C;
    defparam rom3.INIT_RAM_25 = 288'h8743A1D0E85210000000000000000001AD189349A6D369B4DA4D0A854626D46A34DA6D26;
    defparam rom3.INIT_RAM_26 = 288'h8C42A150A8542A150A7E389ACD6A351A8C000035A3D1E8D45A29148A45229148A45A311C;
    defparam rom3.INIT_RAM_27 = 288'h86432190C86000000000000000000000810A8C4DA8D46A351A6D18854626D46A351A8D36;
    defparam rom3.INIT_RAM_28 = 288'h9346231188C462311885389ACD6A351A8C000011A351A8C4622D168B45A2D148A45A311C;
    defparam rom3.INIT_RAM_29 = 288'h8542A21108800000000000000000000000C68549A6D36A351A6D268C49A6D46A351A8D36;
    defparam rom3.INIT_RAM_2A = 288'h9B4DA6D369B4DA6D369B1E8F47A3D1E8F400001122D168C462351A8D46231168A45A311C;
    defparam rom3.INIT_RAM_2B = 288'h8543A25188C00000004139840000000000207342A31269B51A8D369B4DA8D46A351A8D46;
    defparam rom3.INIT_RAM_2C = 288'hA351A8D46A351A8D46A31E8F47A3D1E8F4000033229148B46A3D1E8E47231168A45A311C;
    defparam rom3.INIT_RAM_2D = 288'h8543A2D1C8E088000073429CC400000000001039A15189B51A8D46A351A8D46A351A8D46;
    defparam rom3.INIT_RAM_2E = 288'hA351A8D46A351A8D46A3378F47A3D1E87800234622D168C46A3D1E8E47231188B462311C;
    defparam rom3.INIT_RAM_2F = 288'h8644225168C3C0400010399F8F04F0D0000000081CD0A934DA6D46A351A8D46A351A8D46;
    defparam rom3.INIT_RAM_30 = 288'hA351A8D46A351A8D46A351A8D460000000227C462351A8D47A391C8E472391A8D46A391C;
    defparam rom3.INIT_RAM_31 = 288'h8843A210E87441D02000000ECE26B358F47A1E00040E6854624D36A351A8D46A351A8D46;
    defparam rom3.INIT_RAM_32 = 288'hA351A8D46A351A8D46A351A8D460000044F88E4723D1E8F472391C8E472391E8F47A391C;
    defparam rom3.INIT_RAM_33 = 288'h8A442190A8542A18E81000000BA6B358F47A3D00000208542A3136A351A8D46A351A8D46;
    defparam rom3.INIT_RAM_34 = 288'hA351A8D46A351A8D46A351A8CA200089F11C8C46A3D1E8F472391C8F47A4120904823D1C;
    defparam rom3.INIT_RAM_35 = 288'h8943A1D0C8642A190E7608000186B358F47A1E00000008542A3136A351A8D46A351A8D46;
    defparam rom3.INIT_RAM_36 = 288'h0000000000000000000000000000035239188B462351C8E472391E9149249249248A411E;
    defparam rom3.INIT_RAM_37 = 288'h874421D108743A190E893C040000000000000000000006342A3136A35194400000000000;
    defparam rom3.INIT_RAM_38 = 288'h0000000000000000000000000002347231168A45A311C8E472391E9249A4D2693492411E;
    defparam rom3.INIT_RAM_39 = 288'h8643A25148943A190E89451E0440000000000000000002042A3136A35180000000000000;
    defparam rom3.INIT_RAM_3A = 288'h000000000000000000000000000684622D168A45A351C8E472391E9149249249248A411E;
    defparam rom3.INIT_RAM_3B = 288'h8744225148943A190E8844A25106410800000000000000031A15269B5194400000000000;
    defparam rom3.INIT_RAM_3C = 288'hA351A8D46A351A8D465100000008844225128A45A351E8F472391C904824120904823D1E;
    defparam rom3.INIT_RAM_3D = 288'h8944A29148943A190C8743A1D0E8643A25148B462388E00081CD0A8C49A8D46A351A8D46;
    defparam rom3.INIT_RAM_3E = 288'hA351A8D46A351A8D46A30000020864321D128A45A351E8F472391C8F47A3D1E8F47A3D1E;
    defparam rom3.INIT_RAM_3F = 288'h8A45229148943A190C86432190C8643A25148B462391C0000040C6854626D46A351A8D46;
`endif // _img3_vh_
