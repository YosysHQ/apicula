../img-rom2.vh