`ifndef _img2_vh_
`define _img2_vh_
    defparam rom2.INIT_RAM_00 = 288'h7E3E9F0F87C3F201048341A1104803F201068542209028242215067F3E9F90081412110A;
    defparam rom2.INIT_RAM_01 = 288'h4825138A0552F990CE6C371C0E6753A9E0F27A3D9F4F87D3E9F4FA7C3D9E4F07A3F204FE;
    defparam rom2.INIT_RAM_02 = 288'h7D3E1F0D60038209088341A09048040205088542209028242215067F3E9F90081412110A;
    defparam rom2.INIT_RAM_03 = 288'h4A2593CA0542F188C869361B4E0713A1E0F67B3E1F0FA7E3F9FCFC5C0F000000010180FC;
    defparam rom2.INIT_RAM_04 = 288'h6B3E1AC1E00081CD0A8441205028140A09088542209028242215067F3E9F90081412110A;
    defparam rom2.INIT_RAM_05 = 288'h4B2613CA0542E184C668359B0DC6F391E0F87C3E1F0FA7F409C04000000000000000003C;
    defparam rom2.INIT_RAM_06 = 288'h0F3E03C000000040E682401FCFE7F3FA0104834120D048341A1104803F1FD028241A110A;
    defparam rom2.INIT_RAM_07 = 288'h4A259349E532D984C668359ACDA6E389D4F0783D1E8F67E3803C00000000000000000000;
    defparam rom2.INIT_RAM_08 = 288'h00000003EFF0F80020703F1F4FA7D3E9F4FC7F40A09088341A090480402050684422150A;
    defparam rom2.INIT_RAM_09 = 288'h482492C985015000000006974D66C369C4E4733A9D8EE6B078001862313FDFEFF5F8FC00;
    defparam rom2.INIT_RAM_0A = 288'h1F0007DBEFF6F87C000F359F0F87C3E1F0FA7D3FA0D0A8441205028140A09088542A150C;
    defparam rom2.INIT_RAM_0B = 288'h4724128964B00000000000034A06B361B8DE70399D0AC0E00030AA62313FDFEFF7FBFD7E;
    defparam rom2.INIT_RAM_0C = 288'hDF0037DFEFF7FB7C3E00079ACFC7E3F1F8FC7F40A0D0A844120502824120D088542A150C;
    defparam rom2.INIT_RAM_0D = 288'h4824924944A00000000000000001A289B8DE702A870000006154C47575BFDFEFF7FBFDFE;
    defparam rom2.INIT_RAM_0E = 288'hFF7FBFDFEFF7FBFD7E0000079008241209068341A150A84412050483422110A8542A150C;
    defparam rom2.INIT_RAM_0F = 288'h4A2492490480000000453C044000000000000000000000C2A988C4D77FBFDFEFF7FBFDFE;
    defparam rom2.INIT_RAM_10 = 288'hFF7FBFDFEFF7FBFDFE3F00000C68542A150A8542A150C8541205048442A150A8542A150C;
    defparam rom2.INIT_RAM_11 = 288'h4B251208E47040000078451E000000000000000000030553118910FF7FBFDFEFF7FBFDFE;
    defparam rom2.INIT_RAM_12 = 288'hFF7FBFDFEFF7FBFDFEBF00000428341A0D068341A150A8441A090683422110884422110A;
    defparam rom2.INIT_RAM_13 = 288'h4A2492490471E82000113C2288A000000000001119CEC6C31189AEFF7FBFDFEFF7FBFDFE;
    defparam rom2.INIT_RAM_14 = 288'h7F001FDFEFF7FBFDFEFF00000005F3F9FCFE7F40A0D0A854221106834120904824120904;
    defparam rom2.INIT_RAM_15 = 288'h48249249449238F4100000115148A45229148A45228FE6C31189FEFF7F9FC007F7FBFDFE;
    defparam rom2.INIT_RAM_16 = 288'h0000001FEFF7FBFDFEFF00000001F3E9F4FA7D3FA0D0A8542A15088240A05028140A0502;
    defparam rom2.INIT_RAM_17 = 288'h4724128964A2411C7A0800000F08A45229148A45228FE6C31189FEFF7F80000007FBFDFE;
    defparam rom2.INIT_RAM_18 = 288'h7F001FDFEFF7FBFDFEFF0000000002E9F8FC7E4020D0A8542A15088240A0504824120904;
    defparam rom2.INIT_RAM_19 = 288'h48249249449249208E3D0400022783F9FCFE7F45228FE6C31189FEFF7F9FC007F7FBFDFE;
    defparam rom2.INIT_RAM_1A = 288'hFF7FBFDFEFF7FBFDFED7311881800079BD008040A110A8542A15088240A0906844221108;
    defparam rom2.INIT_RAM_1B = 288'h4A2492490492492892471E8200011339B0D8763FA28FE6C31189AEFF7FBFDFEFF7FBFDFE;
    defparam rom2.INIT_RAM_1C = 288'hFF7FBFDFEFF7FBFDFE8831188AA0C0003CE081412150C86432190A8240A09088542A150A;
    defparam rom2.INIT_RAM_1D = 288'h4B251208E482512C9448238F4100006154C46C3FA28FE6C3118910FF7FBFDFEFF7FBFDFE;
    defparam rom2.INIT_RAM_1E = 288'hFF7FBFDFEFF7FBFDAE62311B0D867088001E70412150C8642A1506834120D088542A150A;
    defparam rom2.INIT_RAM_1F = 288'h4A2492490492512C9449241207E0900030AA623B1FCEC7636188C4D77FBFDFEFF7FBFDFE;
    defparam rom2.INIT_RAM_20 = 288'hEB313ADFEFF7FBACEA623B1FCFE7F3C044000F39A150C8541A09068342A150A8542A150A;
    defparam rom2.INIT_RAM_21 = 288'h4824924944A2592C964A251289441048001855311B0EC763F9D8C47575BFDFEFF7FBFDFE;
    defparam rom2.INIT_RAM_22 = 288'h75311D5D6FF759D4C46C3FA29148A451E02200081D10C85412050485432190C86432190C;
    defparam rom2.INIT_RAM_23 = 288'h4724128964B2592C964B2592C964B20824000C2A988D87F451FCD8623AB5DFEFF7FBFDAE;
    defparam rom2.INIT_RAM_24 = 288'h6231188EAFF3A988D8763B1FCFE7F3FA28F01100040E88541205048342A150A8542A150A;
    defparam rom2.INIT_RAM_25 = 288'h4824924944A2592C964A25128964B250FC100006154D87F451FCEC6C361D94EE16BA20C4;
    defparam rom2.INIT_RAM_26 = 288'h6231188C462311D8FE763B1B0D86C361D9147808800207341205028241209048241A110A;
    defparam rom2.INIT_RAM_27 = 288'h4A2492490492512C944924124944B25120680000060EC7F45228FE7F3F9FD147F36188C4;
    defparam rom2.INIT_RAM_28 = 288'h6231188C462361FD147F36188C462311B0FE8A3C000000F38205028140A050281412110A;
    defparam rom2.INIT_RAM_29 = 288'h4B251208E482512C944823920944B251208E1100000CE8A45229148A45229147F36188C4;
    defparam rom2.INIT_RAM_2A = 288'h6C361B0D86C3B1D8FE7631188C462311B0FE8A451140000079C1048241209048241A110A;
    defparam rom2.INIT_RAM_2B = 288'h4E26928924A25930964924124944B25124903500000448A45229148A3F9FCFE763B1B0D8;
    defparam rom2.INIT_RAM_2C = 288'h7F3F9FCFE7F3B1D8D86218800000000000000022A28F0110003CE48442211088542A150A;
    defparam rom2.INIT_RAM_2D = 288'h54291409C4E2793C9A4B25128964B25928944A00000008A452288A11339B0D8763B1FCFE;
    defparam rom2.INIT_RAM_2E = 288'h8A45229148A3F9B0C462000000000000000000001E1147800000208542A150A86432190C;
    defparam rom2.INIT_RAM_2F = 288'h582B148A050281409E4C2592C964B2592C964B00000008A45228220006154C46C3FA2914;
    defparam rom2.INIT_RAM_30 = 288'h7F3F9FCFE7F3B1B0C46200000000000000000000044F04500000008542A150A86432150A;
    defparam rom2.INIT_RAM_31 = 288'h5C2D164AE572A954A85328944A050281389C4E00000008A45228000000030AA623B1FCFE;
    defparam rom2.INIT_RAM_32 = 288'h6C361B0D86C36188C46200000003E3E9FCC22100000000000000008542A150C8642A150A;
    defparam rom2.INIT_RAM_33 = 288'h6633190C86331180C05F2F978B85B2C95CA85400000008A4522990C80C0001855311B0D8;
    defparam rom2.INIT_RAM_34 = 288'h6231188C46231188C46200000007D3E9FD0685318400000000000086432190C8642A150A;
    defparam rom2.INIT_RAM_35 = 288'h6B359ACD66A33998CC6633190C4612F168B05800000008A4522990C857000000C24988C4;
    defparam rom2.INIT_RAM_36 = 288'h6231188C46231188C46200000007C3E1F90685429D02000000008485432190A854221108;
    defparam rom2.INIT_RAM_37 = 288'h6D369B4DA6C359A8D4683419CCA643117CB85C00000008A4522990C86418C00000006092;
    defparam rom2.INIT_RAM_38 = 288'hC86432000000032190C8000003A793C9F5048542A150C8542A150A854321506824120904;
    defparam rom2.INIT_RAM_39 = 288'h72391C8E472389C4DE6E369B4D66B3519CCC660D000006745228000031B215C180000000;
    defparam rom2.INIT_RAM_3A = 288'hC86432000000032190C800000B2783C1ED0486432190C8542A150A8543215048140A0502;
    defparam rom2.INIT_RAM_3B = 288'h743A1D0E8743A1D0E670379BCDE6F371B0D66B280000022452280000002B990AE0000000;
    defparam rom2.INIT_RAM_3C = 288'h636418C00000018D906300064DE733C1ED048542A150A854221108854321506824120904;
    defparam rom2.INIT_RAM_3D = 288'h753A9D4EA753B1D8EA74391C8E070379B8DA6D38070000033A288A00000615C630000000;
    defparam rom2.INIT_RAM_3E = 288'h0000000000000000000000130D4733C1ED048542A150A8441A090685432150884422110A;
    defparam rom2.INIT_RAM_3F = 288'h773B9DCEE783C9ECF6793C9DCEA73399C8E4723915800000011514780880000000000000;
`endif // _img2_vh_
