`define R_MSB 3
`define G_MSB 3
`define B_MSB 3

