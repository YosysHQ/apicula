`ifndef _img_ram_vh_
`define _img_ram_vh_
    defparam mem.INIT_RAM_00 = 256'h0F0F0F0F0F0F101010101010100F101010101010101010100F0F0F1010101010;
    defparam mem.INIT_RAM_01 = 256'h0909090A0A0B0C0C0D0D0E0E0E0E0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F0F100F;
    defparam mem.INIT_RAM_02 = 256'h0F0F0F0D000E1010101010101010101010101010101010100F0F0F1010101010;
    defparam mem.INIT_RAM_03 = 256'h0909090A0A0B0C0C0D0D0D0E0E0E0F0F0F0F0F0F0F0F0F0F0B03000000040C0F;
    defparam mem.INIT_RAM_04 = 256'h0D0F0D0100020E10101010101010101010101010101010100F0F0F1010101010;
    defparam mem.INIT_RAM_05 = 256'h0909090A0A0B0C0C0D0D0D0D0D0E0F0F0F0F0F0F0F100E040000000000000003;
    defparam mem.INIT_RAM_06 = 256'h010F01000000020E10100F0F0F0F10101010101010101010100F0F1010101010;
    defparam mem.INIT_RAM_07 = 256'h090909090A0B0C0C0D0D0D0D0D0E0E0F0F0F0F0F0F0E01000000000000000000;
    defparam mem.INIT_RAM_08 = 256'h000000031F0300020E0F0F0F0F0F0F0F0F101010101010101010101010101010;
    defparam mem.INIT_RAM_09 = 256'h090909090A05000000010B0D0D0D0E0E0E0E0E0E0D0100010C0C1F1F1F170700;
    defparam mem.INIT_RAM_0A = 256'h0300031B1F1B0300010D0F0F0F0F0F0F0F0F1010101010101010101010101010;
    defparam mem.INIT_RAM_0B = 256'h08090909090000000000010A0D0D0D0D0E0E0E0A0100010A0C0C1F1F1F1F1F17;
    defparam mem.INIT_RAM_0C = 256'h1B001B1F1F1F1B0300010D0F0F0F0F0F0F101010101010101010101010101010;
    defparam mem.INIT_RAM_0D = 256'h090909090900000000000000030A0D0D0E0A030000010A0C0E1D1F1F1F1F1F1F;
    defparam mem.INIT_RAM_0E = 256'h1F1F1F1F1F1F1F17000003101010101010101010101010101010101010101010;
    defparam mem.INIT_RAM_0F = 256'h0909090909000000080F02000000000000000000010A0C0C1A1F1F1F1F1F1F1F;
    defparam mem.INIT_RAM_10 = 256'h1F1F1F1F1F1F1F1F0700000C1010101010101010101010101010101010101010;
    defparam mem.INIT_RAM_11 = 256'h09090908080100000F110F0000000000000000030A0C0C111F1F1F1F1F1F1F1F;
    defparam mem.INIT_RAM_12 = 256'h1F1F1F1F1F1F1F1F170000041010101010101010101010101010101010101010;
    defparam mem.INIT_RAM_13 = 256'h0909090908070100020F11080000000000040C0E0D0C0C1A1F1F1F1F1F1F1F1F;
    defparam mem.INIT_RAM_14 = 256'h0F000F1F1F1F1F1F1F0000000B0F0F0F0F101010101010101010101010101010;
    defparam mem.INIT_RAM_15 = 256'h090909090908070100000811111111111111110F0D0C0C1F1F1F0F000F1F1F1F;
    defparam mem.INIT_RAM_16 = 256'h0000001F1F1F1F1F1F000000030F0F0F0F0F1010101010101010101010101010;
    defparam mem.INIT_RAM_17 = 256'h08090909090908070100000F111111111111110F0D0C0C1F1F1F0000001F1F1F;
    defparam mem.INIT_RAM_18 = 256'h0F000F1F1F1F1F1F1F000000000B0F0F0F101010101010101010101010101010;
    defparam mem.INIT_RAM_19 = 256'h0909090909090908070100020F0F0F0F0F11110F0D0C0C1F1F1F0F000F1F1F1F;
    defparam mem.INIT_RAM_1A = 256'h1F1F1F1F1F1F1F1F1A0C0C0100010D1010101010101010101010101010101010;
    defparam mem.INIT_RAM_1B = 256'h090909090909090908070100020C0D0D0E0F110F0D0C0C1A1F1F1F1F1F1F1F1F;
    defparam mem.INIT_RAM_1C = 256'h1F1F1F1F1F1F1F1F110C0C0A0100010E10101010101010101010101010101010;
    defparam mem.INIT_RAM_1D = 256'h09090908090909090908070100010A0C0D0F110F0D0C0C111F1F1F1F1F1F1F1F;
    defparam mem.INIT_RAM_1E = 256'h1F1F1F1F1F1F1F1A0C0C0D0D0C0200010E101010101010101010101010101010;
    defparam mem.INIT_RAM_1F = 256'h0909090909090909090909070100010A0C0E0F0E0E0D0C0C1A1F1F1F1F1F1F1F;
    defparam mem.INIT_RAM_20 = 256'h1D0C1D1F1F1F1D0E0C0E0F0F0F0F0200010E1010101010101010101010101010;
    defparam mem.INIT_RAM_21 = 256'h090909090909090909090909080100010A0C0D0E0E0F0E0C0E1D1F1F1F1F1F1F;
    defparam mem.INIT_RAM_22 = 256'h0E0C0E1D1F1D0E0C0D0F111111110F0200020E10101010101010101010101010;
    defparam mem.INIT_RAM_23 = 256'h08090909090909090909090909080100010A0C0D0F110F0D0C0E1A1F1F1F1F1A;
    defparam mem.INIT_RAM_24 = 256'h0C0C0C0E1F0E0C0D0E0E0F0F0F0F110F0200020E101010101010101010101010;
    defparam mem.INIT_RAM_25 = 256'h0909090909090909090909090909070100010A0D0F110F0E0D0D0E141C1A110C;
    defparam mem.INIT_RAM_26 = 256'h0C0C0C0C0C0C0E0F0E0E0D0D0D0D0E110F0200020E1010101010101010101010;
    defparam mem.INIT_RAM_27 = 256'h090909090909090909090909090909060000030E0F11110F0F0F0F110F0D0C0C;
    defparam mem.INIT_RAM_28 = 256'h0C0C0C0C0C0D0F110F0D0C0C0C0C0D0F110F0000010E10101010101010101010;
    defparam mem.INIT_RAM_29 = 256'h090909080909090909080909090909080200000C11111111111111110F0D0C0C;
    defparam mem.INIT_RAM_2A = 256'h0D0D0D0D0D0E0E0F0E0C0C0C0C0C0D0F1111080000010E101010101010101010;
    defparam mem.INIT_RAM_2B = 256'h090909090909090909090909090909090600000411111111110F0F0F0E0E0D0D;
    defparam mem.INIT_RAM_2C = 256'h0F0F0F0F0F0E0E0D0C060000000000000008110F0200010E1010101010101010;
    defparam mem.INIT_RAM_2D = 256'h0A0A0A090909090909090909090909090900000011111108020C0D0D0E0E0F0F;
    defparam mem.INIT_RAM_2E = 256'h11111111110F0D0C0C0000000000000000000F110F0000021010101010101010;
    defparam mem.INIT_RAM_2F = 256'h0B0A0A0A0A0A0A090909090909090909090000001111110200010A0C0D0F1111;
    defparam mem.INIT_RAM_30 = 256'h0F0F0F0F0F0E0D0C0C000000000000000000020F080000001010101010101010;
    defparam mem.INIT_RAM_31 = 256'h0B0B0B0A0A0A0A0A0A0A0A0A0A0A090909000000111111000000010A0C0E0F0F;
    defparam mem.INIT_RAM_32 = 256'h0D0D0D0D0D0D0C0C0C000000070F0F0C04000000000000001010101010101010;
    defparam mem.INIT_RAM_33 = 256'h0C0C0C0C0C0C0C0C0B0B0B0B0B0B0A0A0A00000011111119190300010A0C0D0D;
    defparam mem.INIT_RAM_34 = 256'h0C0C0C0C0C0C0C0C0C0000000F0F0F10100C0200000000001010101010101010;
    defparam mem.INIT_RAM_35 = 256'h0D0D0D0D0D0C0C0C0C0C0C0C0C0B0B0B0B000000111111191915000001090C0C;
    defparam mem.INIT_RAM_36 = 256'h0C0C0C0C0C0C0C0C0C0000000F0F0F1010100E02000000081010101010101010;
    defparam mem.INIT_RAM_37 = 256'h0D0D0D0D0D0D0D0D0D0D0C0C0C0C0B0B0B0000001111111919190C0000000309;
    defparam mem.INIT_RAM_38 = 256'h1919190000001919190000030F0F0F1010101010101010101010101010101010;
    defparam mem.INIT_RAM_39 = 256'h0E0E0E0E0E0E0E0D0D0D0D0D0D0D0C0C0C0300000C111100000C191503000000;
    defparam mem.INIT_RAM_3A = 256'h19191900000019191900000B0F0F0F1010101010101010101010101010101010;
    defparam mem.INIT_RAM_3B = 256'h0E0E0E0E0E0E0E0E0E0D0D0D0D0D0D0D0D0A0000041111000000151915000000;
    defparam mem.INIT_RAM_3C = 256'h0C190C0000000C190C00030D0E0F0F1010101010101010101010101010101010;
    defparam mem.INIT_RAM_3D = 256'h0E0E0E0E0E0E0E0E0E0E0E0E0E0D0D0D0D0E0300000C1108000003150C000000;
    defparam mem.INIT_RAM_3E = 256'h00000000000000000000090D0E0F0F1010101010101010101010101010101010;
    defparam mem.INIT_RAM_3F = 256'h0E0E0E0E0F0F0F0F0F0F0E0E0E0E0E0E0E0E0A00000008110F02000000000000;
`endif // _img_ram_h_
