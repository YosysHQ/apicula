module top(O0);
    output O0;
    wire I0;
        OBUF obuf(
            .O(O0),
            .I(I0)
        );
endmodule
// vim: set et ts=4 sw=4:
