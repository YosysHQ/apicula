`define PLL_DYN
`define PLL_DEVICE "GW1N-4"
`define PLL_FCLKIN "12"
`define PLL_ODIV_SEL  64

`define PLL_FBDIV_SEL 12
`define PLL_IDIV_SEL  5

`define PLL_FBDIV_SEL_1 9
`define PLL_IDIV_SEL_1  2

// LCD
`define PLL_FBDIV_SEL_LCD 1
`define PLL_IDIV_SEL_LCD  2

// two pll outputs
`define PLL_0_CLKOUT  PLL_0_CLKOUT 
`define PLL_0_CLKOUTD PLL_0_CLKOUTD
`define PLL_0_LOCK    PLL_0_LOCK   
`define PLL_1_CLKOUT  PLL_1_CLKOUT 
`define PLL_1_CLKOUTD PLL_1_CLKOUTD
`define PLL_1_LOCK    PLL_1_LOCK   
