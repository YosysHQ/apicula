`define R_MSB 4
`define G_MSB 5
`define B_MSB 4

