`define PLL_DYN
`define PLL_DEVICE "GW1NZ-1"
`define PLL_FCLKIN "27"
`define PLL_ODIV_SEL  64

`define PLL_FBDIV_SEL 15
`define PLL_IDIV_SEL  7

`define PLL_FBDIV_SEL_1 0
`define PLL_IDIV_SEL_1  2

// LCD
`define PLL_FBDIV_SEL_LCD 0
`define PLL_IDIV_SEL_LCD  2

