../img-rom3.vh