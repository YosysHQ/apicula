`define PLL_DEVICE "GW1NZ-1"
`define PLL_FCLKIN "27"
`define PLL_FBDIV_SEL 12 // 58.5 MHz (12, 5, 8)  63 MHz (6, 2, 8)
`define PLL_IDIV_SEL  5
`define PLL_ODIV_SEL  8

