`define PLL_DYN
`define PLL_DEVICE "GW1N-1"
`define PLL_FCLKIN "24"
`define PLL_ODIV_SEL  8

`define PLL_FBDIV_SEL 12
`define PLL_IDIV_SEL  5

`define PLL_FBDIV_SEL_1 9
`define PLL_IDIV_SEL_1  2

`define PLL_FBDIV_SEL_LCD 29
`define PLL_IDIV_SEL_LCD   7
