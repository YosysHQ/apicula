../img-rom1.vh